//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9 (64-bit)
//Part Number: GW5AST-LV138PG484AC2/I1
//Device: GW5AST-138B
//Device Version: B
//Created Time: Mon Nov 11 00:57:35 2024

module Gowin_RAM16S (dout, wre, ad, di, clk);

output [2:0] dout;
input wre;
input [13:0] ad;
input [2:0] di;
input clk;

wire ad4_inv;
wire ad5_inv;
wire ad6_inv;
wire lut_f_0;
wire ad7_inv;
wire ad8_inv;
wire ad9_inv;
wire ad10_inv;
wire lut_f_1;
wire ad11_inv;
wire ad12_inv;
wire ad13_inv;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire lut_f_32;
wire lut_f_33;
wire lut_f_34;
wire lut_f_35;
wire lut_f_36;
wire lut_f_37;
wire lut_f_38;
wire lut_f_39;
wire lut_f_40;
wire lut_f_41;
wire lut_f_42;
wire lut_f_43;
wire lut_f_44;
wire lut_f_45;
wire lut_f_46;
wire lut_f_47;
wire lut_f_48;
wire lut_f_49;
wire lut_f_50;
wire lut_f_51;
wire lut_f_52;
wire lut_f_53;
wire lut_f_54;
wire lut_f_55;
wire lut_f_56;
wire lut_f_57;
wire lut_f_58;
wire lut_f_59;
wire lut_f_60;
wire lut_f_61;
wire lut_f_62;
wire lut_f_63;
wire lut_f_64;
wire lut_f_65;
wire lut_f_66;
wire lut_f_67;
wire lut_f_68;
wire lut_f_69;
wire lut_f_70;
wire lut_f_71;
wire lut_f_72;
wire lut_f_73;
wire lut_f_74;
wire lut_f_75;
wire lut_f_76;
wire lut_f_77;
wire lut_f_78;
wire lut_f_79;
wire lut_f_80;
wire lut_f_81;
wire lut_f_82;
wire lut_f_83;
wire lut_f_84;
wire lut_f_85;
wire lut_f_86;
wire lut_f_87;
wire lut_f_88;
wire lut_f_89;
wire lut_f_90;
wire lut_f_91;
wire lut_f_92;
wire lut_f_93;
wire lut_f_94;
wire lut_f_95;
wire lut_f_96;
wire lut_f_97;
wire lut_f_98;
wire lut_f_99;
wire lut_f_100;
wire lut_f_101;
wire lut_f_102;
wire lut_f_103;
wire lut_f_104;
wire lut_f_105;
wire lut_f_106;
wire lut_f_107;
wire lut_f_108;
wire lut_f_109;
wire lut_f_110;
wire lut_f_111;
wire lut_f_112;
wire lut_f_113;
wire lut_f_114;
wire lut_f_115;
wire lut_f_116;
wire lut_f_117;
wire lut_f_118;
wire lut_f_119;
wire lut_f_120;
wire lut_f_121;
wire lut_f_122;
wire lut_f_123;
wire lut_f_124;
wire lut_f_125;
wire lut_f_126;
wire lut_f_127;
wire lut_f_128;
wire lut_f_129;
wire lut_f_130;
wire lut_f_131;
wire lut_f_132;
wire lut_f_133;
wire lut_f_134;
wire lut_f_135;
wire lut_f_136;
wire lut_f_137;
wire lut_f_138;
wire lut_f_139;
wire lut_f_140;
wire lut_f_141;
wire lut_f_142;
wire lut_f_143;
wire lut_f_144;
wire lut_f_145;
wire lut_f_146;
wire lut_f_147;
wire lut_f_148;
wire lut_f_149;
wire lut_f_150;
wire lut_f_151;
wire lut_f_152;
wire lut_f_153;
wire lut_f_154;
wire lut_f_155;
wire lut_f_156;
wire lut_f_157;
wire lut_f_158;
wire lut_f_159;
wire lut_f_160;
wire lut_f_161;
wire lut_f_162;
wire lut_f_163;
wire lut_f_164;
wire lut_f_165;
wire lut_f_166;
wire lut_f_167;
wire lut_f_168;
wire lut_f_169;
wire lut_f_170;
wire lut_f_171;
wire lut_f_172;
wire lut_f_173;
wire lut_f_174;
wire lut_f_175;
wire lut_f_176;
wire lut_f_177;
wire lut_f_178;
wire lut_f_179;
wire lut_f_180;
wire lut_f_181;
wire lut_f_182;
wire lut_f_183;
wire lut_f_184;
wire lut_f_185;
wire lut_f_186;
wire lut_f_187;
wire lut_f_188;
wire lut_f_189;
wire lut_f_190;
wire lut_f_191;
wire lut_f_192;
wire lut_f_193;
wire lut_f_194;
wire lut_f_195;
wire lut_f_196;
wire lut_f_197;
wire lut_f_198;
wire lut_f_199;
wire lut_f_200;
wire lut_f_201;
wire lut_f_202;
wire lut_f_203;
wire lut_f_204;
wire lut_f_205;
wire lut_f_206;
wire lut_f_207;
wire lut_f_208;
wire lut_f_209;
wire lut_f_210;
wire lut_f_211;
wire lut_f_212;
wire lut_f_213;
wire lut_f_214;
wire lut_f_215;
wire lut_f_216;
wire lut_f_217;
wire lut_f_218;
wire lut_f_219;
wire lut_f_220;
wire lut_f_221;
wire lut_f_222;
wire lut_f_223;
wire lut_f_224;
wire lut_f_225;
wire lut_f_226;
wire lut_f_227;
wire lut_f_228;
wire lut_f_229;
wire lut_f_230;
wire lut_f_231;
wire lut_f_232;
wire lut_f_233;
wire lut_f_234;
wire lut_f_235;
wire lut_f_236;
wire lut_f_237;
wire lut_f_238;
wire lut_f_239;
wire lut_f_240;
wire lut_f_241;
wire lut_f_242;
wire lut_f_243;
wire lut_f_244;
wire lut_f_245;
wire lut_f_246;
wire lut_f_247;
wire lut_f_248;
wire lut_f_249;
wire lut_f_250;
wire lut_f_251;
wire lut_f_252;
wire lut_f_253;
wire lut_f_254;
wire lut_f_255;
wire lut_f_256;
wire lut_f_257;
wire lut_f_258;
wire lut_f_259;
wire lut_f_260;
wire lut_f_261;
wire lut_f_262;
wire lut_f_263;
wire lut_f_264;
wire lut_f_265;
wire lut_f_266;
wire lut_f_267;
wire lut_f_268;
wire lut_f_269;
wire lut_f_270;
wire lut_f_271;
wire lut_f_272;
wire lut_f_273;
wire lut_f_274;
wire lut_f_275;
wire lut_f_276;
wire lut_f_277;
wire lut_f_278;
wire lut_f_279;
wire lut_f_280;
wire lut_f_281;
wire lut_f_282;
wire lut_f_283;
wire lut_f_284;
wire lut_f_285;
wire lut_f_286;
wire lut_f_287;
wire lut_f_288;
wire lut_f_289;
wire lut_f_290;
wire lut_f_291;
wire lut_f_292;
wire lut_f_293;
wire lut_f_294;
wire lut_f_295;
wire lut_f_296;
wire lut_f_297;
wire lut_f_298;
wire lut_f_299;
wire lut_f_300;
wire lut_f_301;
wire lut_f_302;
wire lut_f_303;
wire lut_f_304;
wire lut_f_305;
wire lut_f_306;
wire lut_f_307;
wire lut_f_308;
wire lut_f_309;
wire lut_f_310;
wire lut_f_311;
wire lut_f_312;
wire lut_f_313;
wire lut_f_314;
wire lut_f_315;
wire lut_f_316;
wire lut_f_317;
wire lut_f_318;
wire lut_f_319;
wire lut_f_320;
wire lut_f_321;
wire lut_f_322;
wire lut_f_323;
wire lut_f_324;
wire lut_f_325;
wire lut_f_326;
wire lut_f_327;
wire lut_f_328;
wire lut_f_329;
wire lut_f_330;
wire lut_f_331;
wire lut_f_332;
wire lut_f_333;
wire lut_f_334;
wire lut_f_335;
wire lut_f_336;
wire lut_f_337;
wire lut_f_338;
wire lut_f_339;
wire lut_f_340;
wire lut_f_341;
wire lut_f_342;
wire lut_f_343;
wire lut_f_344;
wire lut_f_345;
wire lut_f_346;
wire lut_f_347;
wire lut_f_348;
wire lut_f_349;
wire lut_f_350;
wire lut_f_351;
wire lut_f_352;
wire lut_f_353;
wire lut_f_354;
wire lut_f_355;
wire lut_f_356;
wire lut_f_357;
wire lut_f_358;
wire lut_f_359;
wire lut_f_360;
wire lut_f_361;
wire lut_f_362;
wire lut_f_363;
wire lut_f_364;
wire lut_f_365;
wire lut_f_366;
wire lut_f_367;
wire lut_f_368;
wire lut_f_369;
wire lut_f_370;
wire lut_f_371;
wire lut_f_372;
wire lut_f_373;
wire lut_f_374;
wire lut_f_375;
wire lut_f_376;
wire lut_f_377;
wire lut_f_378;
wire lut_f_379;
wire lut_f_380;
wire lut_f_381;
wire lut_f_382;
wire lut_f_383;
wire lut_f_384;
wire lut_f_385;
wire lut_f_386;
wire lut_f_387;
wire lut_f_388;
wire lut_f_389;
wire lut_f_390;
wire lut_f_391;
wire lut_f_392;
wire lut_f_393;
wire lut_f_394;
wire lut_f_395;
wire lut_f_396;
wire lut_f_397;
wire lut_f_398;
wire lut_f_399;
wire lut_f_400;
wire lut_f_401;
wire lut_f_402;
wire lut_f_403;
wire lut_f_404;
wire lut_f_405;
wire lut_f_406;
wire lut_f_407;
wire lut_f_408;
wire lut_f_409;
wire lut_f_410;
wire lut_f_411;
wire lut_f_412;
wire lut_f_413;
wire lut_f_414;
wire lut_f_415;
wire lut_f_416;
wire lut_f_417;
wire lut_f_418;
wire lut_f_419;
wire lut_f_420;
wire lut_f_421;
wire lut_f_422;
wire lut_f_423;
wire lut_f_424;
wire lut_f_425;
wire lut_f_426;
wire lut_f_427;
wire lut_f_428;
wire lut_f_429;
wire lut_f_430;
wire lut_f_431;
wire lut_f_432;
wire lut_f_433;
wire lut_f_434;
wire lut_f_435;
wire lut_f_436;
wire lut_f_437;
wire lut_f_438;
wire lut_f_439;
wire lut_f_440;
wire lut_f_441;
wire lut_f_442;
wire lut_f_443;
wire lut_f_444;
wire lut_f_445;
wire lut_f_446;
wire lut_f_447;
wire lut_f_448;
wire lut_f_449;
wire lut_f_450;
wire lut_f_451;
wire lut_f_452;
wire lut_f_453;
wire lut_f_454;
wire lut_f_455;
wire lut_f_456;
wire lut_f_457;
wire lut_f_458;
wire lut_f_459;
wire lut_f_460;
wire lut_f_461;
wire lut_f_462;
wire lut_f_463;
wire lut_f_464;
wire lut_f_465;
wire lut_f_466;
wire lut_f_467;
wire lut_f_468;
wire lut_f_469;
wire lut_f_470;
wire lut_f_471;
wire lut_f_472;
wire lut_f_473;
wire lut_f_474;
wire lut_f_475;
wire lut_f_476;
wire lut_f_477;
wire lut_f_478;
wire lut_f_479;
wire lut_f_480;
wire lut_f_481;
wire lut_f_482;
wire lut_f_483;
wire lut_f_484;
wire lut_f_485;
wire lut_f_486;
wire lut_f_487;
wire lut_f_488;
wire lut_f_489;
wire lut_f_490;
wire lut_f_491;
wire lut_f_492;
wire lut_f_493;
wire lut_f_494;
wire lut_f_495;
wire lut_f_496;
wire lut_f_497;
wire lut_f_498;
wire lut_f_499;
wire lut_f_500;
wire lut_f_501;
wire lut_f_502;
wire lut_f_503;
wire lut_f_504;
wire lut_f_505;
wire lut_f_506;
wire lut_f_507;
wire lut_f_508;
wire lut_f_509;
wire lut_f_510;
wire lut_f_511;
wire lut_f_512;
wire lut_f_513;
wire lut_f_514;
wire lut_f_515;
wire lut_f_516;
wire lut_f_517;
wire lut_f_518;
wire lut_f_519;
wire lut_f_520;
wire lut_f_521;
wire lut_f_522;
wire lut_f_523;
wire lut_f_524;
wire lut_f_525;
wire lut_f_526;
wire lut_f_527;
wire lut_f_528;
wire lut_f_529;
wire lut_f_530;
wire lut_f_531;
wire lut_f_532;
wire lut_f_533;
wire lut_f_534;
wire lut_f_535;
wire lut_f_536;
wire lut_f_537;
wire lut_f_538;
wire lut_f_539;
wire lut_f_540;
wire lut_f_541;
wire lut_f_542;
wire lut_f_543;
wire lut_f_544;
wire lut_f_545;
wire lut_f_546;
wire lut_f_547;
wire lut_f_548;
wire lut_f_549;
wire lut_f_550;
wire lut_f_551;
wire lut_f_552;
wire lut_f_553;
wire lut_f_554;
wire lut_f_555;
wire lut_f_556;
wire lut_f_557;
wire lut_f_558;
wire lut_f_559;
wire lut_f_560;
wire lut_f_561;
wire lut_f_562;
wire lut_f_563;
wire lut_f_564;
wire lut_f_565;
wire lut_f_566;
wire lut_f_567;
wire lut_f_568;
wire lut_f_569;
wire lut_f_570;
wire lut_f_571;
wire lut_f_572;
wire lut_f_573;
wire lut_f_574;
wire lut_f_575;
wire lut_f_576;
wire lut_f_577;
wire lut_f_578;
wire lut_f_579;
wire lut_f_580;
wire lut_f_581;
wire lut_f_582;
wire lut_f_583;
wire lut_f_584;
wire lut_f_585;
wire lut_f_586;
wire lut_f_587;
wire lut_f_588;
wire lut_f_589;
wire lut_f_590;
wire lut_f_591;
wire lut_f_592;
wire lut_f_593;
wire lut_f_594;
wire lut_f_595;
wire lut_f_596;
wire lut_f_597;
wire lut_f_598;
wire lut_f_599;
wire lut_f_600;
wire lut_f_601;
wire lut_f_602;
wire lut_f_603;
wire lut_f_604;
wire lut_f_605;
wire lut_f_606;
wire lut_f_607;
wire lut_f_608;
wire lut_f_609;
wire lut_f_610;
wire lut_f_611;
wire lut_f_612;
wire lut_f_613;
wire lut_f_614;
wire lut_f_615;
wire lut_f_616;
wire lut_f_617;
wire lut_f_618;
wire lut_f_619;
wire lut_f_620;
wire lut_f_621;
wire lut_f_622;
wire lut_f_623;
wire lut_f_624;
wire lut_f_625;
wire lut_f_626;
wire lut_f_627;
wire lut_f_628;
wire lut_f_629;
wire lut_f_630;
wire lut_f_631;
wire lut_f_632;
wire lut_f_633;
wire lut_f_634;
wire lut_f_635;
wire lut_f_636;
wire lut_f_637;
wire lut_f_638;
wire lut_f_639;
wire lut_f_640;
wire lut_f_641;
wire lut_f_642;
wire lut_f_643;
wire lut_f_644;
wire lut_f_645;
wire lut_f_646;
wire lut_f_647;
wire lut_f_648;
wire lut_f_649;
wire lut_f_650;
wire lut_f_651;
wire lut_f_652;
wire lut_f_653;
wire lut_f_654;
wire lut_f_655;
wire lut_f_656;
wire lut_f_657;
wire lut_f_658;
wire lut_f_659;
wire lut_f_660;
wire lut_f_661;
wire lut_f_662;
wire lut_f_663;
wire lut_f_664;
wire lut_f_665;
wire lut_f_666;
wire lut_f_667;
wire lut_f_668;
wire lut_f_669;
wire lut_f_670;
wire lut_f_671;
wire lut_f_672;
wire lut_f_673;
wire lut_f_674;
wire lut_f_675;
wire lut_f_676;
wire lut_f_677;
wire lut_f_678;
wire lut_f_679;
wire lut_f_680;
wire lut_f_681;
wire lut_f_682;
wire lut_f_683;
wire lut_f_684;
wire lut_f_685;
wire lut_f_686;
wire lut_f_687;
wire lut_f_688;
wire lut_f_689;
wire lut_f_690;
wire lut_f_691;
wire lut_f_692;
wire lut_f_693;
wire lut_f_694;
wire lut_f_695;
wire lut_f_696;
wire lut_f_697;
wire lut_f_698;
wire lut_f_699;
wire lut_f_700;
wire lut_f_701;
wire lut_f_702;
wire lut_f_703;
wire lut_f_704;
wire lut_f_705;
wire lut_f_706;
wire lut_f_707;
wire lut_f_708;
wire lut_f_709;
wire lut_f_710;
wire lut_f_711;
wire lut_f_712;
wire lut_f_713;
wire lut_f_714;
wire lut_f_715;
wire lut_f_716;
wire lut_f_717;
wire lut_f_718;
wire lut_f_719;
wire lut_f_720;
wire lut_f_721;
wire lut_f_722;
wire lut_f_723;
wire lut_f_724;
wire lut_f_725;
wire lut_f_726;
wire lut_f_727;
wire lut_f_728;
wire lut_f_729;
wire lut_f_730;
wire lut_f_731;
wire lut_f_732;
wire lut_f_733;
wire lut_f_734;
wire lut_f_735;
wire lut_f_736;
wire lut_f_737;
wire lut_f_738;
wire lut_f_739;
wire lut_f_740;
wire lut_f_741;
wire lut_f_742;
wire lut_f_743;
wire lut_f_744;
wire lut_f_745;
wire lut_f_746;
wire lut_f_747;
wire lut_f_748;
wire lut_f_749;
wire lut_f_750;
wire lut_f_751;
wire lut_f_752;
wire lut_f_753;
wire lut_f_754;
wire lut_f_755;
wire lut_f_756;
wire lut_f_757;
wire lut_f_758;
wire lut_f_759;
wire lut_f_760;
wire lut_f_761;
wire lut_f_762;
wire lut_f_763;
wire lut_f_764;
wire lut_f_765;
wire lut_f_766;
wire lut_f_767;
wire lut_f_768;
wire lut_f_769;
wire lut_f_770;
wire lut_f_771;
wire lut_f_772;
wire lut_f_773;
wire lut_f_774;
wire lut_f_775;
wire lut_f_776;
wire lut_f_777;
wire lut_f_778;
wire lut_f_779;
wire lut_f_780;
wire lut_f_781;
wire lut_f_782;
wire lut_f_783;
wire lut_f_784;
wire lut_f_785;
wire lut_f_786;
wire lut_f_787;
wire lut_f_788;
wire lut_f_789;
wire lut_f_790;
wire lut_f_791;
wire lut_f_792;
wire lut_f_793;
wire lut_f_794;
wire lut_f_795;
wire lut_f_796;
wire lut_f_797;
wire lut_f_798;
wire lut_f_799;
wire lut_f_800;
wire lut_f_801;
wire lut_f_802;
wire lut_f_803;
wire lut_f_804;
wire lut_f_805;
wire lut_f_806;
wire lut_f_807;
wire lut_f_808;
wire lut_f_809;
wire lut_f_810;
wire lut_f_811;
wire lut_f_812;
wire lut_f_813;
wire lut_f_814;
wire lut_f_815;
wire lut_f_816;
wire lut_f_817;
wire lut_f_818;
wire lut_f_819;
wire lut_f_820;
wire lut_f_821;
wire lut_f_822;
wire lut_f_823;
wire lut_f_824;
wire lut_f_825;
wire lut_f_826;
wire lut_f_827;
wire lut_f_828;
wire lut_f_829;
wire lut_f_830;
wire lut_f_831;
wire lut_f_832;
wire lut_f_833;
wire lut_f_834;
wire lut_f_835;
wire lut_f_836;
wire lut_f_837;
wire lut_f_838;
wire lut_f_839;
wire lut_f_840;
wire lut_f_841;
wire lut_f_842;
wire lut_f_843;
wire lut_f_844;
wire lut_f_845;
wire lut_f_846;
wire lut_f_847;
wire lut_f_848;
wire lut_f_849;
wire lut_f_850;
wire lut_f_851;
wire lut_f_852;
wire lut_f_853;
wire lut_f_854;
wire lut_f_855;
wire lut_f_856;
wire lut_f_857;
wire lut_f_858;
wire lut_f_859;
wire lut_f_860;
wire lut_f_861;
wire lut_f_862;
wire lut_f_863;
wire lut_f_864;
wire lut_f_865;
wire lut_f_866;
wire lut_f_867;
wire lut_f_868;
wire lut_f_869;
wire lut_f_870;
wire lut_f_871;
wire lut_f_872;
wire lut_f_873;
wire lut_f_874;
wire lut_f_875;
wire lut_f_876;
wire lut_f_877;
wire lut_f_878;
wire lut_f_879;
wire lut_f_880;
wire lut_f_881;
wire lut_f_882;
wire lut_f_883;
wire lut_f_884;
wire lut_f_885;
wire lut_f_886;
wire lut_f_887;
wire lut_f_888;
wire lut_f_889;
wire lut_f_890;
wire lut_f_891;
wire lut_f_892;
wire lut_f_893;
wire lut_f_894;
wire lut_f_895;
wire lut_f_896;
wire lut_f_897;
wire lut_f_898;
wire lut_f_899;
wire lut_f_900;
wire lut_f_901;
wire lut_f_902;
wire lut_f_903;
wire lut_f_904;
wire lut_f_905;
wire lut_f_906;
wire lut_f_907;
wire lut_f_908;
wire lut_f_909;
wire lut_f_910;
wire lut_f_911;
wire lut_f_912;
wire lut_f_913;
wire lut_f_914;
wire lut_f_915;
wire lut_f_916;
wire lut_f_917;
wire lut_f_918;
wire lut_f_919;
wire lut_f_920;
wire lut_f_921;
wire lut_f_922;
wire lut_f_923;
wire lut_f_924;
wire lut_f_925;
wire lut_f_926;
wire lut_f_927;
wire lut_f_928;
wire lut_f_929;
wire lut_f_930;
wire lut_f_931;
wire lut_f_932;
wire lut_f_933;
wire lut_f_934;
wire lut_f_935;
wire lut_f_936;
wire lut_f_937;
wire lut_f_938;
wire lut_f_939;
wire lut_f_940;
wire lut_f_941;
wire lut_f_942;
wire lut_f_943;
wire lut_f_944;
wire lut_f_945;
wire lut_f_946;
wire lut_f_947;
wire lut_f_948;
wire lut_f_949;
wire lut_f_950;
wire lut_f_951;
wire lut_f_952;
wire lut_f_953;
wire lut_f_954;
wire lut_f_955;
wire lut_f_956;
wire lut_f_957;
wire lut_f_958;
wire lut_f_959;
wire lut_f_960;
wire lut_f_961;
wire lut_f_962;
wire lut_f_963;
wire lut_f_964;
wire lut_f_965;
wire lut_f_966;
wire lut_f_967;
wire lut_f_968;
wire lut_f_969;
wire lut_f_970;
wire lut_f_971;
wire lut_f_972;
wire lut_f_973;
wire lut_f_974;
wire lut_f_975;
wire lut_f_976;
wire lut_f_977;
wire lut_f_978;
wire lut_f_979;
wire lut_f_980;
wire lut_f_981;
wire lut_f_982;
wire lut_f_983;
wire lut_f_984;
wire lut_f_985;
wire lut_f_986;
wire lut_f_987;
wire lut_f_988;
wire lut_f_989;
wire lut_f_990;
wire lut_f_991;
wire lut_f_992;
wire lut_f_993;
wire lut_f_994;
wire lut_f_995;
wire lut_f_996;
wire lut_f_997;
wire lut_f_998;
wire lut_f_999;
wire lut_f_1000;
wire lut_f_1001;
wire lut_f_1002;
wire lut_f_1003;
wire lut_f_1004;
wire lut_f_1005;
wire lut_f_1006;
wire lut_f_1007;
wire lut_f_1008;
wire lut_f_1009;
wire lut_f_1010;
wire lut_f_1011;
wire lut_f_1012;
wire lut_f_1013;
wire lut_f_1014;
wire lut_f_1015;
wire lut_f_1016;
wire lut_f_1017;
wire lut_f_1018;
wire lut_f_1019;
wire lut_f_1020;
wire lut_f_1021;
wire lut_f_1022;
wire lut_f_1023;
wire lut_f_1024;
wire lut_f_1025;
wire lut_f_1026;
wire lut_f_1027;
wire lut_f_1028;
wire lut_f_1029;
wire lut_f_1030;
wire lut_f_1031;
wire lut_f_1032;
wire lut_f_1033;
wire lut_f_1034;
wire lut_f_1035;
wire lut_f_1036;
wire lut_f_1037;
wire lut_f_1038;
wire lut_f_1039;
wire lut_f_1040;
wire lut_f_1041;
wire lut_f_1042;
wire lut_f_1043;
wire lut_f_1044;
wire lut_f_1045;
wire lut_f_1046;
wire lut_f_1047;
wire lut_f_1048;
wire lut_f_1049;
wire lut_f_1050;
wire lut_f_1051;
wire lut_f_1052;
wire lut_f_1053;
wire lut_f_1054;
wire lut_f_1055;
wire lut_f_1056;
wire lut_f_1057;
wire lut_f_1058;
wire lut_f_1059;
wire lut_f_1060;
wire lut_f_1061;
wire lut_f_1062;
wire lut_f_1063;
wire lut_f_1064;
wire lut_f_1065;
wire lut_f_1066;
wire lut_f_1067;
wire lut_f_1068;
wire lut_f_1069;
wire lut_f_1070;
wire lut_f_1071;
wire lut_f_1072;
wire lut_f_1073;
wire lut_f_1074;
wire lut_f_1075;
wire lut_f_1076;
wire lut_f_1077;
wire lut_f_1078;
wire lut_f_1079;
wire lut_f_1080;
wire lut_f_1081;
wire lut_f_1082;
wire lut_f_1083;
wire lut_f_1084;
wire lut_f_1085;
wire lut_f_1086;
wire lut_f_1087;
wire lut_f_1088;
wire lut_f_1089;
wire lut_f_1090;
wire lut_f_1091;
wire lut_f_1092;
wire lut_f_1093;
wire lut_f_1094;
wire lut_f_1095;
wire lut_f_1096;
wire lut_f_1097;
wire lut_f_1098;
wire lut_f_1099;
wire lut_f_1100;
wire lut_f_1101;
wire lut_f_1102;
wire lut_f_1103;
wire lut_f_1104;
wire lut_f_1105;
wire lut_f_1106;
wire lut_f_1107;
wire lut_f_1108;
wire lut_f_1109;
wire lut_f_1110;
wire lut_f_1111;
wire lut_f_1112;
wire lut_f_1113;
wire lut_f_1114;
wire lut_f_1115;
wire lut_f_1116;
wire lut_f_1117;
wire lut_f_1118;
wire lut_f_1119;
wire lut_f_1120;
wire lut_f_1121;
wire lut_f_1122;
wire lut_f_1123;
wire lut_f_1124;
wire lut_f_1125;
wire lut_f_1126;
wire lut_f_1127;
wire lut_f_1128;
wire lut_f_1129;
wire lut_f_1130;
wire lut_f_1131;
wire lut_f_1132;
wire lut_f_1133;
wire lut_f_1134;
wire lut_f_1135;
wire lut_f_1136;
wire lut_f_1137;
wire lut_f_1138;
wire lut_f_1139;
wire lut_f_1140;
wire lut_f_1141;
wire lut_f_1142;
wire lut_f_1143;
wire lut_f_1144;
wire lut_f_1145;
wire lut_f_1146;
wire lut_f_1147;
wire lut_f_1148;
wire lut_f_1149;
wire lut_f_1150;
wire lut_f_1151;
wire lut_f_1152;
wire lut_f_1153;
wire lut_f_1154;
wire lut_f_1155;
wire lut_f_1156;
wire lut_f_1157;
wire lut_f_1158;
wire lut_f_1159;
wire lut_f_1160;
wire lut_f_1161;
wire lut_f_1162;
wire lut_f_1163;
wire lut_f_1164;
wire lut_f_1165;
wire lut_f_1166;
wire lut_f_1167;
wire lut_f_1168;
wire lut_f_1169;
wire lut_f_1170;
wire lut_f_1171;
wire lut_f_1172;
wire lut_f_1173;
wire lut_f_1174;
wire lut_f_1175;
wire lut_f_1176;
wire lut_f_1177;
wire lut_f_1178;
wire lut_f_1179;
wire lut_f_1180;
wire lut_f_1181;
wire lut_f_1182;
wire lut_f_1183;
wire lut_f_1184;
wire lut_f_1185;
wire lut_f_1186;
wire lut_f_1187;
wire lut_f_1188;
wire lut_f_1189;
wire lut_f_1190;
wire lut_f_1191;
wire lut_f_1192;
wire lut_f_1193;
wire lut_f_1194;
wire lut_f_1195;
wire lut_f_1196;
wire lut_f_1197;
wire lut_f_1198;
wire lut_f_1199;
wire lut_f_1200;
wire lut_f_1201;
wire lut_f_1202;
wire lut_f_1203;
wire lut_f_1204;
wire lut_f_1205;
wire lut_f_1206;
wire lut_f_1207;
wire lut_f_1208;
wire lut_f_1209;
wire lut_f_1210;
wire lut_f_1211;
wire lut_f_1212;
wire lut_f_1213;
wire lut_f_1214;
wire lut_f_1215;
wire lut_f_1216;
wire lut_f_1217;
wire lut_f_1218;
wire lut_f_1219;
wire lut_f_1220;
wire lut_f_1221;
wire lut_f_1222;
wire lut_f_1223;
wire lut_f_1224;
wire lut_f_1225;
wire lut_f_1226;
wire lut_f_1227;
wire lut_f_1228;
wire lut_f_1229;
wire lut_f_1230;
wire lut_f_1231;
wire lut_f_1232;
wire lut_f_1233;
wire lut_f_1234;
wire lut_f_1235;
wire lut_f_1236;
wire lut_f_1237;
wire lut_f_1238;
wire lut_f_1239;
wire lut_f_1240;
wire lut_f_1241;
wire lut_f_1242;
wire lut_f_1243;
wire lut_f_1244;
wire lut_f_1245;
wire lut_f_1246;
wire lut_f_1247;
wire lut_f_1248;
wire lut_f_1249;
wire lut_f_1250;
wire lut_f_1251;
wire lut_f_1252;
wire lut_f_1253;
wire lut_f_1254;
wire lut_f_1255;
wire lut_f_1256;
wire lut_f_1257;
wire lut_f_1258;
wire lut_f_1259;
wire lut_f_1260;
wire lut_f_1261;
wire lut_f_1262;
wire lut_f_1263;
wire lut_f_1264;
wire lut_f_1265;
wire lut_f_1266;
wire lut_f_1267;
wire lut_f_1268;
wire lut_f_1269;
wire lut_f_1270;
wire lut_f_1271;
wire lut_f_1272;
wire lut_f_1273;
wire lut_f_1274;
wire lut_f_1275;
wire lut_f_1276;
wire lut_f_1277;
wire lut_f_1278;
wire lut_f_1279;
wire lut_f_1280;
wire lut_f_1281;
wire lut_f_1282;
wire lut_f_1283;
wire lut_f_1284;
wire lut_f_1285;
wire lut_f_1286;
wire lut_f_1287;
wire lut_f_1288;
wire lut_f_1289;
wire lut_f_1290;
wire lut_f_1291;
wire lut_f_1292;
wire lut_f_1293;
wire lut_f_1294;
wire lut_f_1295;
wire lut_f_1296;
wire lut_f_1297;
wire lut_f_1298;
wire lut_f_1299;
wire lut_f_1300;
wire lut_f_1301;
wire lut_f_1302;
wire lut_f_1303;
wire lut_f_1304;
wire lut_f_1305;
wire lut_f_1306;
wire lut_f_1307;
wire lut_f_1308;
wire lut_f_1309;
wire lut_f_1310;
wire lut_f_1311;
wire lut_f_1312;
wire lut_f_1313;
wire lut_f_1314;
wire lut_f_1315;
wire lut_f_1316;
wire lut_f_1317;
wire lut_f_1318;
wire lut_f_1319;
wire lut_f_1320;
wire lut_f_1321;
wire lut_f_1322;
wire lut_f_1323;
wire lut_f_1324;
wire lut_f_1325;
wire lut_f_1326;
wire lut_f_1327;
wire lut_f_1328;
wire lut_f_1329;
wire lut_f_1330;
wire lut_f_1331;
wire lut_f_1332;
wire lut_f_1333;
wire lut_f_1334;
wire lut_f_1335;
wire lut_f_1336;
wire lut_f_1337;
wire lut_f_1338;
wire lut_f_1339;
wire lut_f_1340;
wire lut_f_1341;
wire lut_f_1342;
wire lut_f_1343;
wire lut_f_1344;
wire lut_f_1345;
wire lut_f_1346;
wire lut_f_1347;
wire lut_f_1348;
wire lut_f_1349;
wire lut_f_1350;
wire lut_f_1351;
wire lut_f_1352;
wire lut_f_1353;
wire lut_f_1354;
wire lut_f_1355;
wire lut_f_1356;
wire lut_f_1357;
wire lut_f_1358;
wire lut_f_1359;
wire lut_f_1360;
wire lut_f_1361;
wire lut_f_1362;
wire lut_f_1363;
wire lut_f_1364;
wire lut_f_1365;
wire lut_f_1366;
wire lut_f_1367;
wire lut_f_1368;
wire lut_f_1369;
wire lut_f_1370;
wire lut_f_1371;
wire lut_f_1372;
wire lut_f_1373;
wire lut_f_1374;
wire lut_f_1375;
wire lut_f_1376;
wire lut_f_1377;
wire lut_f_1378;
wire lut_f_1379;
wire lut_f_1380;
wire lut_f_1381;
wire lut_f_1382;
wire lut_f_1383;
wire lut_f_1384;
wire lut_f_1385;
wire lut_f_1386;
wire lut_f_1387;
wire lut_f_1388;
wire lut_f_1389;
wire lut_f_1390;
wire lut_f_1391;
wire lut_f_1392;
wire lut_f_1393;
wire lut_f_1394;
wire lut_f_1395;
wire lut_f_1396;
wire lut_f_1397;
wire lut_f_1398;
wire lut_f_1399;
wire lut_f_1400;
wire lut_f_1401;
wire lut_f_1402;
wire lut_f_1403;
wire lut_f_1404;
wire lut_f_1405;
wire lut_f_1406;
wire lut_f_1407;
wire lut_f_1408;
wire lut_f_1409;
wire lut_f_1410;
wire lut_f_1411;
wire lut_f_1412;
wire lut_f_1413;
wire lut_f_1414;
wire lut_f_1415;
wire lut_f_1416;
wire lut_f_1417;
wire lut_f_1418;
wire lut_f_1419;
wire lut_f_1420;
wire lut_f_1421;
wire lut_f_1422;
wire lut_f_1423;
wire lut_f_1424;
wire lut_f_1425;
wire lut_f_1426;
wire lut_f_1427;
wire lut_f_1428;
wire lut_f_1429;
wire lut_f_1430;
wire lut_f_1431;
wire lut_f_1432;
wire lut_f_1433;
wire lut_f_1434;
wire lut_f_1435;
wire lut_f_1436;
wire lut_f_1437;
wire lut_f_1438;
wire lut_f_1439;
wire lut_f_1440;
wire lut_f_1441;
wire lut_f_1442;
wire lut_f_1443;
wire lut_f_1444;
wire lut_f_1445;
wire lut_f_1446;
wire lut_f_1447;
wire lut_f_1448;
wire lut_f_1449;
wire lut_f_1450;
wire lut_f_1451;
wire lut_f_1452;
wire lut_f_1453;
wire lut_f_1454;
wire lut_f_1455;
wire lut_f_1456;
wire lut_f_1457;
wire lut_f_1458;
wire lut_f_1459;
wire lut_f_1460;
wire lut_f_1461;
wire lut_f_1462;
wire lut_f_1463;
wire lut_f_1464;
wire lut_f_1465;
wire lut_f_1466;
wire lut_f_1467;
wire lut_f_1468;
wire lut_f_1469;
wire lut_f_1470;
wire lut_f_1471;
wire lut_f_1472;
wire lut_f_1473;
wire lut_f_1474;
wire lut_f_1475;
wire lut_f_1476;
wire lut_f_1477;
wire lut_f_1478;
wire lut_f_1479;
wire lut_f_1480;
wire lut_f_1481;
wire lut_f_1482;
wire lut_f_1483;
wire lut_f_1484;
wire lut_f_1485;
wire lut_f_1486;
wire lut_f_1487;
wire lut_f_1488;
wire lut_f_1489;
wire lut_f_1490;
wire lut_f_1491;
wire lut_f_1492;
wire lut_f_1493;
wire lut_f_1494;
wire lut_f_1495;
wire lut_f_1496;
wire lut_f_1497;
wire lut_f_1498;
wire lut_f_1499;
wire lut_f_1500;
wire lut_f_1501;
wire lut_f_1502;
wire lut_f_1503;
wire lut_f_1504;
wire lut_f_1505;
wire lut_f_1506;
wire lut_f_1507;
wire lut_f_1508;
wire lut_f_1509;
wire lut_f_1510;
wire lut_f_1511;
wire lut_f_1512;
wire lut_f_1513;
wire lut_f_1514;
wire lut_f_1515;
wire lut_f_1516;
wire lut_f_1517;
wire lut_f_1518;
wire lut_f_1519;
wire lut_f_1520;
wire lut_f_1521;
wire lut_f_1522;
wire lut_f_1523;
wire lut_f_1524;
wire lut_f_1525;
wire lut_f_1526;
wire lut_f_1527;
wire lut_f_1528;
wire lut_f_1529;
wire lut_f_1530;
wire lut_f_1531;
wire lut_f_1532;
wire lut_f_1533;
wire lut_f_1534;
wire lut_f_1535;
wire lut_f_1536;
wire lut_f_1537;
wire lut_f_1538;
wire lut_f_1539;
wire lut_f_1540;
wire lut_f_1541;
wire lut_f_1542;
wire lut_f_1543;
wire lut_f_1544;
wire lut_f_1545;
wire lut_f_1546;
wire lut_f_1547;
wire lut_f_1548;
wire lut_f_1549;
wire lut_f_1550;
wire lut_f_1551;
wire lut_f_1552;
wire lut_f_1553;
wire lut_f_1554;
wire lut_f_1555;
wire lut_f_1556;
wire lut_f_1557;
wire lut_f_1558;
wire lut_f_1559;
wire lut_f_1560;
wire lut_f_1561;
wire lut_f_1562;
wire lut_f_1563;
wire lut_f_1564;
wire lut_f_1565;
wire lut_f_1566;
wire lut_f_1567;
wire lut_f_1568;
wire lut_f_1569;
wire lut_f_1570;
wire lut_f_1571;
wire lut_f_1572;
wire lut_f_1573;
wire lut_f_1574;
wire lut_f_1575;
wire lut_f_1576;
wire lut_f_1577;
wire lut_f_1578;
wire lut_f_1579;
wire lut_f_1580;
wire lut_f_1581;
wire lut_f_1582;
wire lut_f_1583;
wire lut_f_1584;
wire lut_f_1585;
wire lut_f_1586;
wire lut_f_1587;
wire lut_f_1588;
wire lut_f_1589;
wire lut_f_1590;
wire lut_f_1591;
wire lut_f_1592;
wire lut_f_1593;
wire lut_f_1594;
wire lut_f_1595;
wire lut_f_1596;
wire lut_f_1597;
wire lut_f_1598;
wire lut_f_1599;
wire lut_f_1600;
wire lut_f_1601;
wire lut_f_1602;
wire lut_f_1603;
wire lut_f_1604;
wire lut_f_1605;
wire lut_f_1606;
wire lut_f_1607;
wire lut_f_1608;
wire lut_f_1609;
wire lut_f_1610;
wire lut_f_1611;
wire lut_f_1612;
wire lut_f_1613;
wire lut_f_1614;
wire lut_f_1615;
wire lut_f_1616;
wire lut_f_1617;
wire lut_f_1618;
wire lut_f_1619;
wire lut_f_1620;
wire lut_f_1621;
wire lut_f_1622;
wire lut_f_1623;
wire lut_f_1624;
wire lut_f_1625;
wire lut_f_1626;
wire lut_f_1627;
wire lut_f_1628;
wire lut_f_1629;
wire lut_f_1630;
wire lut_f_1631;
wire lut_f_1632;
wire lut_f_1633;
wire lut_f_1634;
wire lut_f_1635;
wire lut_f_1636;
wire lut_f_1637;
wire lut_f_1638;
wire lut_f_1639;
wire lut_f_1640;
wire lut_f_1641;
wire lut_f_1642;
wire lut_f_1643;
wire lut_f_1644;
wire lut_f_1645;
wire lut_f_1646;
wire lut_f_1647;
wire lut_f_1648;
wire lut_f_1649;
wire lut_f_1650;
wire lut_f_1651;
wire lut_f_1652;
wire lut_f_1653;
wire lut_f_1654;
wire lut_f_1655;
wire lut_f_1656;
wire lut_f_1657;
wire lut_f_1658;
wire lut_f_1659;
wire lut_f_1660;
wire lut_f_1661;
wire lut_f_1662;
wire lut_f_1663;
wire lut_f_1664;
wire lut_f_1665;
wire lut_f_1666;
wire lut_f_1667;
wire lut_f_1668;
wire lut_f_1669;
wire lut_f_1670;
wire lut_f_1671;
wire lut_f_1672;
wire lut_f_1673;
wire lut_f_1674;
wire lut_f_1675;
wire lut_f_1676;
wire lut_f_1677;
wire lut_f_1678;
wire lut_f_1679;
wire lut_f_1680;
wire lut_f_1681;
wire lut_f_1682;
wire lut_f_1683;
wire lut_f_1684;
wire lut_f_1685;
wire lut_f_1686;
wire lut_f_1687;
wire lut_f_1688;
wire lut_f_1689;
wire lut_f_1690;
wire lut_f_1691;
wire lut_f_1692;
wire lut_f_1693;
wire lut_f_1694;
wire lut_f_1695;
wire lut_f_1696;
wire lut_f_1697;
wire lut_f_1698;
wire lut_f_1699;
wire lut_f_1700;
wire lut_f_1701;
wire lut_f_1702;
wire lut_f_1703;
wire lut_f_1704;
wire lut_f_1705;
wire lut_f_1706;
wire lut_f_1707;
wire lut_f_1708;
wire lut_f_1709;
wire lut_f_1710;
wire lut_f_1711;
wire lut_f_1712;
wire lut_f_1713;
wire lut_f_1714;
wire lut_f_1715;
wire lut_f_1716;
wire lut_f_1717;
wire lut_f_1718;
wire lut_f_1719;
wire lut_f_1720;
wire lut_f_1721;
wire lut_f_1722;
wire lut_f_1723;
wire lut_f_1724;
wire lut_f_1725;
wire lut_f_1726;
wire lut_f_1727;
wire lut_f_1728;
wire lut_f_1729;
wire lut_f_1730;
wire lut_f_1731;
wire lut_f_1732;
wire lut_f_1733;
wire lut_f_1734;
wire lut_f_1735;
wire lut_f_1736;
wire lut_f_1737;
wire lut_f_1738;
wire lut_f_1739;
wire lut_f_1740;
wire lut_f_1741;
wire lut_f_1742;
wire lut_f_1743;
wire lut_f_1744;
wire lut_f_1745;
wire lut_f_1746;
wire lut_f_1747;
wire lut_f_1748;
wire lut_f_1749;
wire lut_f_1750;
wire lut_f_1751;
wire lut_f_1752;
wire lut_f_1753;
wire lut_f_1754;
wire lut_f_1755;
wire lut_f_1756;
wire lut_f_1757;
wire lut_f_1758;
wire lut_f_1759;
wire lut_f_1760;
wire lut_f_1761;
wire lut_f_1762;
wire lut_f_1763;
wire lut_f_1764;
wire lut_f_1765;
wire lut_f_1766;
wire lut_f_1767;
wire lut_f_1768;
wire lut_f_1769;
wire lut_f_1770;
wire lut_f_1771;
wire lut_f_1772;
wire lut_f_1773;
wire lut_f_1774;
wire lut_f_1775;
wire lut_f_1776;
wire lut_f_1777;
wire lut_f_1778;
wire lut_f_1779;
wire lut_f_1780;
wire lut_f_1781;
wire lut_f_1782;
wire lut_f_1783;
wire lut_f_1784;
wire lut_f_1785;
wire lut_f_1786;
wire lut_f_1787;
wire lut_f_1788;
wire lut_f_1789;
wire lut_f_1790;
wire lut_f_1791;
wire lut_f_1792;
wire lut_f_1793;
wire lut_f_1794;
wire lut_f_1795;
wire lut_f_1796;
wire lut_f_1797;
wire lut_f_1798;
wire lut_f_1799;
wire lut_f_1800;
wire lut_f_1801;
wire lut_f_1802;
wire lut_f_1803;
wire lut_f_1804;
wire lut_f_1805;
wire lut_f_1806;
wire lut_f_1807;
wire lut_f_1808;
wire lut_f_1809;
wire lut_f_1810;
wire lut_f_1811;
wire lut_f_1812;
wire lut_f_1813;
wire lut_f_1814;
wire lut_f_1815;
wire lut_f_1816;
wire lut_f_1817;
wire lut_f_1818;
wire lut_f_1819;
wire lut_f_1820;
wire lut_f_1821;
wire lut_f_1822;
wire lut_f_1823;
wire lut_f_1824;
wire lut_f_1825;
wire lut_f_1826;
wire lut_f_1827;
wire lut_f_1828;
wire lut_f_1829;
wire lut_f_1830;
wire lut_f_1831;
wire lut_f_1832;
wire lut_f_1833;
wire lut_f_1834;
wire lut_f_1835;
wire lut_f_1836;
wire lut_f_1837;
wire lut_f_1838;
wire lut_f_1839;
wire lut_f_1840;
wire lut_f_1841;
wire lut_f_1842;
wire lut_f_1843;
wire lut_f_1844;
wire lut_f_1845;
wire lut_f_1846;
wire lut_f_1847;
wire lut_f_1848;
wire lut_f_1849;
wire lut_f_1850;
wire lut_f_1851;
wire lut_f_1852;
wire lut_f_1853;
wire lut_f_1854;
wire lut_f_1855;
wire lut_f_1856;
wire lut_f_1857;
wire lut_f_1858;
wire lut_f_1859;
wire lut_f_1860;
wire lut_f_1861;
wire lut_f_1862;
wire lut_f_1863;
wire lut_f_1864;
wire lut_f_1865;
wire lut_f_1866;
wire lut_f_1867;
wire lut_f_1868;
wire lut_f_1869;
wire lut_f_1870;
wire lut_f_1871;
wire lut_f_1872;
wire lut_f_1873;
wire lut_f_1874;
wire lut_f_1875;
wire lut_f_1876;
wire lut_f_1877;
wire lut_f_1878;
wire lut_f_1879;
wire lut_f_1880;
wire lut_f_1881;
wire lut_f_1882;
wire lut_f_1883;
wire lut_f_1884;
wire lut_f_1885;
wire lut_f_1886;
wire lut_f_1887;
wire lut_f_1888;
wire lut_f_1889;
wire lut_f_1890;
wire lut_f_1891;
wire lut_f_1892;
wire lut_f_1893;
wire lut_f_1894;
wire lut_f_1895;
wire lut_f_1896;
wire lut_f_1897;
wire lut_f_1898;
wire lut_f_1899;
wire lut_f_1900;
wire lut_f_1901;
wire lut_f_1902;
wire lut_f_1903;
wire lut_f_1904;
wire lut_f_1905;
wire lut_f_1906;
wire lut_f_1907;
wire lut_f_1908;
wire lut_f_1909;
wire lut_f_1910;
wire lut_f_1911;
wire lut_f_1912;
wire lut_f_1913;
wire lut_f_1914;
wire lut_f_1915;
wire lut_f_1916;
wire lut_f_1917;
wire lut_f_1918;
wire lut_f_1919;
wire lut_f_1920;
wire lut_f_1921;
wire lut_f_1922;
wire lut_f_1923;
wire lut_f_1924;
wire lut_f_1925;
wire lut_f_1926;
wire lut_f_1927;
wire lut_f_1928;
wire lut_f_1929;
wire lut_f_1930;
wire lut_f_1931;
wire lut_f_1932;
wire lut_f_1933;
wire lut_f_1934;
wire lut_f_1935;
wire lut_f_1936;
wire lut_f_1937;
wire lut_f_1938;
wire lut_f_1939;
wire lut_f_1940;
wire lut_f_1941;
wire lut_f_1942;
wire lut_f_1943;
wire lut_f_1944;
wire lut_f_1945;
wire lut_f_1946;
wire lut_f_1947;
wire lut_f_1948;
wire lut_f_1949;
wire lut_f_1950;
wire lut_f_1951;
wire lut_f_1952;
wire lut_f_1953;
wire lut_f_1954;
wire lut_f_1955;
wire lut_f_1956;
wire lut_f_1957;
wire lut_f_1958;
wire lut_f_1959;
wire lut_f_1960;
wire lut_f_1961;
wire lut_f_1962;
wire lut_f_1963;
wire lut_f_1964;
wire lut_f_1965;
wire lut_f_1966;
wire lut_f_1967;
wire lut_f_1968;
wire lut_f_1969;
wire lut_f_1970;
wire lut_f_1971;
wire lut_f_1972;
wire lut_f_1973;
wire lut_f_1974;
wire lut_f_1975;
wire lut_f_1976;
wire lut_f_1977;
wire lut_f_1978;
wire lut_f_1979;
wire lut_f_1980;
wire lut_f_1981;
wire lut_f_1982;
wire lut_f_1983;
wire lut_f_1984;
wire lut_f_1985;
wire lut_f_1986;
wire lut_f_1987;
wire lut_f_1988;
wire lut_f_1989;
wire lut_f_1990;
wire lut_f_1991;
wire lut_f_1992;
wire lut_f_1993;
wire lut_f_1994;
wire lut_f_1995;
wire lut_f_1996;
wire lut_f_1997;
wire lut_f_1998;
wire lut_f_1999;
wire lut_f_2000;
wire lut_f_2001;
wire lut_f_2002;
wire lut_f_2003;
wire lut_f_2004;
wire lut_f_2005;
wire lut_f_2006;
wire lut_f_2007;
wire lut_f_2008;
wire lut_f_2009;
wire lut_f_2010;
wire lut_f_2011;
wire lut_f_2012;
wire lut_f_2013;
wire lut_f_2014;
wire lut_f_2015;
wire lut_f_2016;
wire lut_f_2017;
wire lut_f_2018;
wire lut_f_2019;
wire lut_f_2020;
wire lut_f_2021;
wire lut_f_2022;
wire lut_f_2023;
wire lut_f_2024;
wire lut_f_2025;
wire lut_f_2026;
wire lut_f_2027;
wire lut_f_2028;
wire lut_f_2029;
wire lut_f_2030;
wire lut_f_2031;
wire lut_f_2032;
wire lut_f_2033;
wire lut_f_2034;
wire lut_f_2035;
wire lut_f_2036;
wire lut_f_2037;
wire lut_f_2038;
wire lut_f_2039;
wire lut_f_2040;
wire lut_f_2041;
wire lut_f_2042;
wire lut_f_2043;
wire lut_f_2044;
wire lut_f_2045;
wire lut_f_2046;
wire lut_f_2047;
wire lut_f_2048;
wire lut_f_2049;
wire lut_f_2050;
wire lut_f_2051;
wire lut_f_2052;
wire lut_f_2053;
wire lut_f_2054;
wire lut_f_2055;
wire lut_f_2056;
wire lut_f_2057;
wire lut_f_2058;
wire lut_f_2059;
wire lut_f_2060;
wire lut_f_2061;
wire lut_f_2062;
wire lut_f_2063;
wire lut_f_2064;
wire lut_f_2065;
wire lut_f_2066;
wire lut_f_2067;
wire lut_f_2068;
wire lut_f_2069;
wire lut_f_2070;
wire lut_f_2071;
wire lut_f_2072;
wire lut_f_2073;
wire lut_f_2074;
wire lut_f_2075;
wire lut_f_2076;
wire lut_f_2077;
wire lut_f_2078;
wire lut_f_2079;
wire lut_f_2080;
wire lut_f_2081;
wire lut_f_2082;
wire lut_f_2083;
wire lut_f_2084;
wire lut_f_2085;
wire lut_f_2086;
wire lut_f_2087;
wire lut_f_2088;
wire lut_f_2089;
wire lut_f_2090;
wire lut_f_2091;
wire lut_f_2092;
wire lut_f_2093;
wire lut_f_2094;
wire lut_f_2095;
wire lut_f_2096;
wire lut_f_2097;
wire lut_f_2098;
wire lut_f_2099;
wire lut_f_2100;
wire lut_f_2101;
wire lut_f_2102;
wire lut_f_2103;
wire lut_f_2104;
wire lut_f_2105;
wire lut_f_2106;
wire lut_f_2107;
wire lut_f_2108;
wire lut_f_2109;
wire lut_f_2110;
wire lut_f_2111;
wire lut_f_2112;
wire lut_f_2113;
wire lut_f_2114;
wire lut_f_2115;
wire lut_f_2116;
wire lut_f_2117;
wire lut_f_2118;
wire lut_f_2119;
wire lut_f_2120;
wire lut_f_2121;
wire lut_f_2122;
wire lut_f_2123;
wire lut_f_2124;
wire lut_f_2125;
wire lut_f_2126;
wire lut_f_2127;
wire lut_f_2128;
wire lut_f_2129;
wire lut_f_2130;
wire lut_f_2131;
wire lut_f_2132;
wire lut_f_2133;
wire lut_f_2134;
wire lut_f_2135;
wire lut_f_2136;
wire lut_f_2137;
wire lut_f_2138;
wire lut_f_2139;
wire lut_f_2140;
wire lut_f_2141;
wire lut_f_2142;
wire lut_f_2143;
wire lut_f_2144;
wire lut_f_2145;
wire lut_f_2146;
wire lut_f_2147;
wire lut_f_2148;
wire lut_f_2149;
wire lut_f_2150;
wire lut_f_2151;
wire lut_f_2152;
wire lut_f_2153;
wire lut_f_2154;
wire lut_f_2155;
wire lut_f_2156;
wire lut_f_2157;
wire lut_f_2158;
wire lut_f_2159;
wire lut_f_2160;
wire lut_f_2161;
wire lut_f_2162;
wire lut_f_2163;
wire lut_f_2164;
wire lut_f_2165;
wire lut_f_2166;
wire lut_f_2167;
wire lut_f_2168;
wire lut_f_2169;
wire lut_f_2170;
wire lut_f_2171;
wire lut_f_2172;
wire lut_f_2173;
wire lut_f_2174;
wire lut_f_2175;
wire lut_f_2176;
wire lut_f_2177;
wire lut_f_2178;
wire lut_f_2179;
wire lut_f_2180;
wire lut_f_2181;
wire lut_f_2182;
wire lut_f_2183;
wire lut_f_2184;
wire lut_f_2185;
wire lut_f_2186;
wire lut_f_2187;
wire lut_f_2188;
wire lut_f_2189;
wire lut_f_2190;
wire lut_f_2191;
wire lut_f_2192;
wire lut_f_2193;
wire lut_f_2194;
wire lut_f_2195;
wire lut_f_2196;
wire lut_f_2197;
wire lut_f_2198;
wire lut_f_2199;
wire lut_f_2200;
wire lut_f_2201;
wire lut_f_2202;
wire lut_f_2203;
wire lut_f_2204;
wire lut_f_2205;
wire lut_f_2206;
wire lut_f_2207;
wire lut_f_2208;
wire lut_f_2209;
wire lut_f_2210;
wire lut_f_2211;
wire lut_f_2212;
wire lut_f_2213;
wire lut_f_2214;
wire lut_f_2215;
wire lut_f_2216;
wire lut_f_2217;
wire lut_f_2218;
wire lut_f_2219;
wire lut_f_2220;
wire lut_f_2221;
wire lut_f_2222;
wire lut_f_2223;
wire lut_f_2224;
wire lut_f_2225;
wire lut_f_2226;
wire lut_f_2227;
wire lut_f_2228;
wire lut_f_2229;
wire lut_f_2230;
wire lut_f_2231;
wire lut_f_2232;
wire lut_f_2233;
wire lut_f_2234;
wire lut_f_2235;
wire lut_f_2236;
wire lut_f_2237;
wire lut_f_2238;
wire lut_f_2239;
wire lut_f_2240;
wire lut_f_2241;
wire lut_f_2242;
wire lut_f_2243;
wire lut_f_2244;
wire lut_f_2245;
wire lut_f_2246;
wire lut_f_2247;
wire lut_f_2248;
wire lut_f_2249;
wire lut_f_2250;
wire lut_f_2251;
wire lut_f_2252;
wire lut_f_2253;
wire lut_f_2254;
wire lut_f_2255;
wire lut_f_2256;
wire lut_f_2257;
wire lut_f_2258;
wire lut_f_2259;
wire lut_f_2260;
wire lut_f_2261;
wire lut_f_2262;
wire lut_f_2263;
wire lut_f_2264;
wire lut_f_2265;
wire lut_f_2266;
wire lut_f_2267;
wire lut_f_2268;
wire lut_f_2269;
wire lut_f_2270;
wire lut_f_2271;
wire lut_f_2272;
wire lut_f_2273;
wire lut_f_2274;
wire lut_f_2275;
wire lut_f_2276;
wire lut_f_2277;
wire lut_f_2278;
wire lut_f_2279;
wire lut_f_2280;
wire lut_f_2281;
wire lut_f_2282;
wire lut_f_2283;
wire lut_f_2284;
wire lut_f_2285;
wire lut_f_2286;
wire lut_f_2287;
wire lut_f_2288;
wire lut_f_2289;
wire lut_f_2290;
wire lut_f_2291;
wire lut_f_2292;
wire lut_f_2293;
wire lut_f_2294;
wire lut_f_2295;
wire lut_f_2296;
wire lut_f_2297;
wire lut_f_2298;
wire lut_f_2299;
wire lut_f_2300;
wire lut_f_2301;
wire lut_f_2302;
wire lut_f_2303;
wire lut_f_2304;
wire lut_f_2305;
wire lut_f_2306;
wire lut_f_2307;
wire lut_f_2308;
wire lut_f_2309;
wire lut_f_2310;
wire lut_f_2311;
wire lut_f_2312;
wire lut_f_2313;
wire lut_f_2314;
wire lut_f_2315;
wire lut_f_2316;
wire lut_f_2317;
wire lut_f_2318;
wire lut_f_2319;
wire lut_f_2320;
wire lut_f_2321;
wire lut_f_2322;
wire lut_f_2323;
wire lut_f_2324;
wire lut_f_2325;
wire lut_f_2326;
wire lut_f_2327;
wire lut_f_2328;
wire lut_f_2329;
wire lut_f_2330;
wire lut_f_2331;
wire lut_f_2332;
wire lut_f_2333;
wire lut_f_2334;
wire lut_f_2335;
wire lut_f_2336;
wire lut_f_2337;
wire lut_f_2338;
wire lut_f_2339;
wire lut_f_2340;
wire lut_f_2341;
wire lut_f_2342;
wire lut_f_2343;
wire lut_f_2344;
wire lut_f_2345;
wire lut_f_2346;
wire lut_f_2347;
wire lut_f_2348;
wire lut_f_2349;
wire lut_f_2350;
wire lut_f_2351;
wire lut_f_2352;
wire lut_f_2353;
wire lut_f_2354;
wire lut_f_2355;
wire lut_f_2356;
wire lut_f_2357;
wire lut_f_2358;
wire lut_f_2359;
wire lut_f_2360;
wire lut_f_2361;
wire lut_f_2362;
wire lut_f_2363;
wire lut_f_2364;
wire lut_f_2365;
wire lut_f_2366;
wire lut_f_2367;
wire lut_f_2368;
wire lut_f_2369;
wire lut_f_2370;
wire lut_f_2371;
wire lut_f_2372;
wire lut_f_2373;
wire lut_f_2374;
wire lut_f_2375;
wire lut_f_2376;
wire lut_f_2377;
wire lut_f_2378;
wire lut_f_2379;
wire lut_f_2380;
wire lut_f_2381;
wire lut_f_2382;
wire lut_f_2383;
wire lut_f_2384;
wire lut_f_2385;
wire lut_f_2386;
wire lut_f_2387;
wire lut_f_2388;
wire lut_f_2389;
wire lut_f_2390;
wire lut_f_2391;
wire lut_f_2392;
wire lut_f_2393;
wire lut_f_2394;
wire lut_f_2395;
wire lut_f_2396;
wire lut_f_2397;
wire lut_f_2398;
wire lut_f_2399;
wire lut_f_2400;
wire lut_f_2401;
wire lut_f_2402;
wire lut_f_2403;
wire lut_f_2404;
wire lut_f_2405;
wire lut_f_2406;
wire lut_f_2407;
wire lut_f_2408;
wire lut_f_2409;
wire lut_f_2410;
wire lut_f_2411;
wire lut_f_2412;
wire lut_f_2413;
wire lut_f_2414;
wire lut_f_2415;
wire lut_f_2416;
wire lut_f_2417;
wire lut_f_2418;
wire lut_f_2419;
wire lut_f_2420;
wire lut_f_2421;
wire lut_f_2422;
wire lut_f_2423;
wire lut_f_2424;
wire lut_f_2425;
wire lut_f_2426;
wire lut_f_2427;
wire lut_f_2428;
wire lut_f_2429;
wire lut_f_2430;
wire lut_f_2431;
wire lut_f_2432;
wire lut_f_2433;
wire lut_f_2434;
wire lut_f_2435;
wire lut_f_2436;
wire lut_f_2437;
wire lut_f_2438;
wire lut_f_2439;
wire lut_f_2440;
wire lut_f_2441;
wire lut_f_2442;
wire lut_f_2443;
wire lut_f_2444;
wire lut_f_2445;
wire lut_f_2446;
wire lut_f_2447;
wire lut_f_2448;
wire lut_f_2449;
wire lut_f_2450;
wire lut_f_2451;
wire lut_f_2452;
wire lut_f_2453;
wire lut_f_2454;
wire lut_f_2455;
wire lut_f_2456;
wire lut_f_2457;
wire lut_f_2458;
wire lut_f_2459;
wire lut_f_2460;
wire lut_f_2461;
wire lut_f_2462;
wire lut_f_2463;
wire lut_f_2464;
wire lut_f_2465;
wire lut_f_2466;
wire lut_f_2467;
wire lut_f_2468;
wire lut_f_2469;
wire lut_f_2470;
wire lut_f_2471;
wire lut_f_2472;
wire lut_f_2473;
wire lut_f_2474;
wire lut_f_2475;
wire lut_f_2476;
wire lut_f_2477;
wire lut_f_2478;
wire lut_f_2479;
wire lut_f_2480;
wire lut_f_2481;
wire lut_f_2482;
wire lut_f_2483;
wire lut_f_2484;
wire lut_f_2485;
wire lut_f_2486;
wire lut_f_2487;
wire lut_f_2488;
wire lut_f_2489;
wire lut_f_2490;
wire lut_f_2491;
wire lut_f_2492;
wire lut_f_2493;
wire lut_f_2494;
wire lut_f_2495;
wire lut_f_2496;
wire lut_f_2497;
wire lut_f_2498;
wire lut_f_2499;
wire lut_f_2500;
wire lut_f_2501;
wire lut_f_2502;
wire lut_f_2503;
wire lut_f_2504;
wire lut_f_2505;
wire lut_f_2506;
wire lut_f_2507;
wire lut_f_2508;
wire lut_f_2509;
wire lut_f_2510;
wire lut_f_2511;
wire lut_f_2512;
wire lut_f_2513;
wire lut_f_2514;
wire lut_f_2515;
wire lut_f_2516;
wire lut_f_2517;
wire lut_f_2518;
wire lut_f_2519;
wire lut_f_2520;
wire lut_f_2521;
wire lut_f_2522;
wire lut_f_2523;
wire lut_f_2524;
wire lut_f_2525;
wire lut_f_2526;
wire lut_f_2527;
wire lut_f_2528;
wire lut_f_2529;
wire lut_f_2530;
wire lut_f_2531;
wire lut_f_2532;
wire lut_f_2533;
wire lut_f_2534;
wire lut_f_2535;
wire lut_f_2536;
wire lut_f_2537;
wire lut_f_2538;
wire lut_f_2539;
wire lut_f_2540;
wire lut_f_2541;
wire lut_f_2542;
wire lut_f_2543;
wire lut_f_2544;
wire lut_f_2545;
wire lut_f_2546;
wire lut_f_2547;
wire lut_f_2548;
wire lut_f_2549;
wire lut_f_2550;
wire lut_f_2551;
wire lut_f_2552;
wire lut_f_2553;
wire lut_f_2554;
wire lut_f_2555;
wire lut_f_2556;
wire lut_f_2557;
wire lut_f_2558;
wire lut_f_2559;
wire lut_f_2560;
wire lut_f_2561;
wire lut_f_2562;
wire lut_f_2563;
wire lut_f_2564;
wire lut_f_2565;
wire lut_f_2566;
wire lut_f_2567;
wire lut_f_2568;
wire lut_f_2569;
wire lut_f_2570;
wire lut_f_2571;
wire lut_f_2572;
wire lut_f_2573;
wire lut_f_2574;
wire lut_f_2575;
wire lut_f_2576;
wire lut_f_2577;
wire lut_f_2578;
wire lut_f_2579;
wire lut_f_2580;
wire lut_f_2581;
wire lut_f_2582;
wire lut_f_2583;
wire lut_f_2584;
wire lut_f_2585;
wire lut_f_2586;
wire lut_f_2587;
wire lut_f_2588;
wire lut_f_2589;
wire lut_f_2590;
wire lut_f_2591;
wire lut_f_2592;
wire lut_f_2593;
wire lut_f_2594;
wire lut_f_2595;
wire lut_f_2596;
wire lut_f_2597;
wire lut_f_2598;
wire lut_f_2599;
wire lut_f_2600;
wire lut_f_2601;
wire lut_f_2602;
wire lut_f_2603;
wire lut_f_2604;
wire lut_f_2605;
wire lut_f_2606;
wire lut_f_2607;
wire lut_f_2608;
wire lut_f_2609;
wire lut_f_2610;
wire lut_f_2611;
wire lut_f_2612;
wire lut_f_2613;
wire lut_f_2614;
wire lut_f_2615;
wire lut_f_2616;
wire lut_f_2617;
wire lut_f_2618;
wire lut_f_2619;
wire lut_f_2620;
wire lut_f_2621;
wire lut_f_2622;
wire lut_f_2623;
wire lut_f_2624;
wire lut_f_2625;
wire lut_f_2626;
wire lut_f_2627;
wire lut_f_2628;
wire lut_f_2629;
wire lut_f_2630;
wire lut_f_2631;
wire lut_f_2632;
wire lut_f_2633;
wire lut_f_2634;
wire lut_f_2635;
wire lut_f_2636;
wire lut_f_2637;
wire lut_f_2638;
wire lut_f_2639;
wire lut_f_2640;
wire lut_f_2641;
wire lut_f_2642;
wire lut_f_2643;
wire lut_f_2644;
wire lut_f_2645;
wire lut_f_2646;
wire lut_f_2647;
wire lut_f_2648;
wire lut_f_2649;
wire lut_f_2650;
wire lut_f_2651;
wire lut_f_2652;
wire lut_f_2653;
wire lut_f_2654;
wire lut_f_2655;
wire lut_f_2656;
wire lut_f_2657;
wire lut_f_2658;
wire lut_f_2659;
wire lut_f_2660;
wire lut_f_2661;
wire lut_f_2662;
wire lut_f_2663;
wire lut_f_2664;
wire lut_f_2665;
wire lut_f_2666;
wire lut_f_2667;
wire lut_f_2668;
wire lut_f_2669;
wire lut_f_2670;
wire lut_f_2671;
wire lut_f_2672;
wire lut_f_2673;
wire lut_f_2674;
wire lut_f_2675;
wire lut_f_2676;
wire lut_f_2677;
wire lut_f_2678;
wire lut_f_2679;
wire lut_f_2680;
wire lut_f_2681;
wire lut_f_2682;
wire lut_f_2683;
wire lut_f_2684;
wire lut_f_2685;
wire lut_f_2686;
wire lut_f_2687;
wire lut_f_2688;
wire lut_f_2689;
wire lut_f_2690;
wire lut_f_2691;
wire lut_f_2692;
wire lut_f_2693;
wire lut_f_2694;
wire lut_f_2695;
wire lut_f_2696;
wire lut_f_2697;
wire lut_f_2698;
wire lut_f_2699;
wire lut_f_2700;
wire lut_f_2701;
wire lut_f_2702;
wire lut_f_2703;
wire lut_f_2704;
wire lut_f_2705;
wire lut_f_2706;
wire lut_f_2707;
wire lut_f_2708;
wire lut_f_2709;
wire lut_f_2710;
wire lut_f_2711;
wire lut_f_2712;
wire lut_f_2713;
wire lut_f_2714;
wire lut_f_2715;
wire lut_f_2716;
wire lut_f_2717;
wire lut_f_2718;
wire lut_f_2719;
wire lut_f_2720;
wire lut_f_2721;
wire lut_f_2722;
wire lut_f_2723;
wire lut_f_2724;
wire lut_f_2725;
wire lut_f_2726;
wire lut_f_2727;
wire lut_f_2728;
wire lut_f_2729;
wire lut_f_2730;
wire lut_f_2731;
wire lut_f_2732;
wire lut_f_2733;
wire lut_f_2734;
wire lut_f_2735;
wire lut_f_2736;
wire lut_f_2737;
wire lut_f_2738;
wire lut_f_2739;
wire lut_f_2740;
wire lut_f_2741;
wire lut_f_2742;
wire lut_f_2743;
wire lut_f_2744;
wire lut_f_2745;
wire lut_f_2746;
wire lut_f_2747;
wire lut_f_2748;
wire lut_f_2749;
wire lut_f_2750;
wire lut_f_2751;
wire lut_f_2752;
wire lut_f_2753;
wire lut_f_2754;
wire lut_f_2755;
wire lut_f_2756;
wire lut_f_2757;
wire lut_f_2758;
wire lut_f_2759;
wire lut_f_2760;
wire lut_f_2761;
wire lut_f_2762;
wire lut_f_2763;
wire lut_f_2764;
wire lut_f_2765;
wire lut_f_2766;
wire lut_f_2767;
wire lut_f_2768;
wire lut_f_2769;
wire lut_f_2770;
wire lut_f_2771;
wire lut_f_2772;
wire lut_f_2773;
wire lut_f_2774;
wire lut_f_2775;
wire lut_f_2776;
wire lut_f_2777;
wire lut_f_2778;
wire lut_f_2779;
wire lut_f_2780;
wire lut_f_2781;
wire lut_f_2782;
wire lut_f_2783;
wire lut_f_2784;
wire lut_f_2785;
wire lut_f_2786;
wire lut_f_2787;
wire lut_f_2788;
wire lut_f_2789;
wire lut_f_2790;
wire lut_f_2791;
wire lut_f_2792;
wire lut_f_2793;
wire lut_f_2794;
wire lut_f_2795;
wire lut_f_2796;
wire lut_f_2797;
wire lut_f_2798;
wire lut_f_2799;
wire lut_f_2800;
wire lut_f_2801;
wire lut_f_2802;
wire lut_f_2803;
wire lut_f_2804;
wire lut_f_2805;
wire lut_f_2806;
wire lut_f_2807;
wire lut_f_2808;
wire lut_f_2809;
wire lut_f_2810;
wire lut_f_2811;
wire lut_f_2812;
wire lut_f_2813;
wire lut_f_2814;
wire lut_f_2815;
wire lut_f_2816;
wire lut_f_2817;
wire lut_f_2818;
wire lut_f_2819;
wire lut_f_2820;
wire lut_f_2821;
wire lut_f_2822;
wire lut_f_2823;
wire lut_f_2824;
wire lut_f_2825;
wire lut_f_2826;
wire lut_f_2827;
wire lut_f_2828;
wire lut_f_2829;
wire lut_f_2830;
wire lut_f_2831;
wire lut_f_2832;
wire lut_f_2833;
wire lut_f_2834;
wire lut_f_2835;
wire lut_f_2836;
wire lut_f_2837;
wire lut_f_2838;
wire lut_f_2839;
wire lut_f_2840;
wire lut_f_2841;
wire lut_f_2842;
wire lut_f_2843;
wire lut_f_2844;
wire lut_f_2845;
wire lut_f_2846;
wire lut_f_2847;
wire lut_f_2848;
wire lut_f_2849;
wire lut_f_2850;
wire lut_f_2851;
wire lut_f_2852;
wire lut_f_2853;
wire lut_f_2854;
wire lut_f_2855;
wire lut_f_2856;
wire lut_f_2857;
wire lut_f_2858;
wire lut_f_2859;
wire lut_f_2860;
wire lut_f_2861;
wire lut_f_2862;
wire lut_f_2863;
wire lut_f_2864;
wire lut_f_2865;
wire lut_f_2866;
wire lut_f_2867;
wire lut_f_2868;
wire lut_f_2869;
wire lut_f_2870;
wire lut_f_2871;
wire lut_f_2872;
wire lut_f_2873;
wire lut_f_2874;
wire lut_f_2875;
wire lut_f_2876;
wire lut_f_2877;
wire lut_f_2878;
wire lut_f_2879;
wire lut_f_2880;
wire lut_f_2881;
wire lut_f_2882;
wire lut_f_2883;
wire lut_f_2884;
wire lut_f_2885;
wire lut_f_2886;
wire lut_f_2887;
wire lut_f_2888;
wire lut_f_2889;
wire lut_f_2890;
wire lut_f_2891;
wire lut_f_2892;
wire lut_f_2893;
wire lut_f_2894;
wire lut_f_2895;
wire lut_f_2896;
wire lut_f_2897;
wire lut_f_2898;
wire lut_f_2899;
wire lut_f_2900;
wire lut_f_2901;
wire lut_f_2902;
wire lut_f_2903;
wire lut_f_2904;
wire lut_f_2905;
wire lut_f_2906;
wire lut_f_2907;
wire lut_f_2908;
wire lut_f_2909;
wire lut_f_2910;
wire lut_f_2911;
wire lut_f_2912;
wire lut_f_2913;
wire lut_f_2914;
wire lut_f_2915;
wire lut_f_2916;
wire lut_f_2917;
wire lut_f_2918;
wire lut_f_2919;
wire lut_f_2920;
wire lut_f_2921;
wire lut_f_2922;
wire lut_f_2923;
wire lut_f_2924;
wire lut_f_2925;
wire lut_f_2926;
wire lut_f_2927;
wire lut_f_2928;
wire lut_f_2929;
wire lut_f_2930;
wire lut_f_2931;
wire lut_f_2932;
wire lut_f_2933;
wire lut_f_2934;
wire lut_f_2935;
wire lut_f_2936;
wire lut_f_2937;
wire lut_f_2938;
wire lut_f_2939;
wire lut_f_2940;
wire lut_f_2941;
wire lut_f_2942;
wire lut_f_2943;
wire lut_f_2944;
wire lut_f_2945;
wire lut_f_2946;
wire lut_f_2947;
wire lut_f_2948;
wire lut_f_2949;
wire lut_f_2950;
wire lut_f_2951;
wire lut_f_2952;
wire lut_f_2953;
wire lut_f_2954;
wire lut_f_2955;
wire lut_f_2956;
wire lut_f_2957;
wire lut_f_2958;
wire lut_f_2959;
wire lut_f_2960;
wire lut_f_2961;
wire lut_f_2962;
wire lut_f_2963;
wire lut_f_2964;
wire lut_f_2965;
wire lut_f_2966;
wire lut_f_2967;
wire lut_f_2968;
wire lut_f_2969;
wire lut_f_2970;
wire lut_f_2971;
wire lut_f_2972;
wire lut_f_2973;
wire lut_f_2974;
wire lut_f_2975;
wire lut_f_2976;
wire lut_f_2977;
wire lut_f_2978;
wire lut_f_2979;
wire lut_f_2980;
wire lut_f_2981;
wire lut_f_2982;
wire lut_f_2983;
wire lut_f_2984;
wire lut_f_2985;
wire lut_f_2986;
wire lut_f_2987;
wire lut_f_2988;
wire lut_f_2989;
wire lut_f_2990;
wire lut_f_2991;
wire lut_f_2992;
wire lut_f_2993;
wire lut_f_2994;
wire lut_f_2995;
wire lut_f_2996;
wire lut_f_2997;
wire lut_f_2998;
wire lut_f_2999;
wire lut_f_3000;
wire lut_f_3001;
wire lut_f_3002;
wire lut_f_3003;
wire lut_f_3004;
wire lut_f_3005;
wire lut_f_3006;
wire lut_f_3007;
wire lut_f_3008;
wire lut_f_3009;
wire lut_f_3010;
wire lut_f_3011;
wire lut_f_3012;
wire lut_f_3013;
wire lut_f_3014;
wire lut_f_3015;
wire lut_f_3016;
wire lut_f_3017;
wire lut_f_3018;
wire lut_f_3019;
wire lut_f_3020;
wire lut_f_3021;
wire lut_f_3022;
wire lut_f_3023;
wire lut_f_3024;
wire lut_f_3025;
wire lut_f_3026;
wire lut_f_3027;
wire lut_f_3028;
wire lut_f_3029;
wire lut_f_3030;
wire lut_f_3031;
wire lut_f_3032;
wire lut_f_3033;
wire lut_f_3034;
wire lut_f_3035;
wire lut_f_3036;
wire lut_f_3037;
wire lut_f_3038;
wire lut_f_3039;
wire lut_f_3040;
wire lut_f_3041;
wire lut_f_3042;
wire lut_f_3043;
wire lut_f_3044;
wire lut_f_3045;
wire lut_f_3046;
wire lut_f_3047;
wire lut_f_3048;
wire lut_f_3049;
wire lut_f_3050;
wire lut_f_3051;
wire lut_f_3052;
wire lut_f_3053;
wire lut_f_3054;
wire lut_f_3055;
wire lut_f_3056;
wire lut_f_3057;
wire lut_f_3058;
wire lut_f_3059;
wire lut_f_3060;
wire lut_f_3061;
wire lut_f_3062;
wire lut_f_3063;
wire lut_f_3064;
wire lut_f_3065;
wire lut_f_3066;
wire lut_f_3067;
wire lut_f_3068;
wire lut_f_3069;
wire lut_f_3070;
wire lut_f_3071;
wire lut_f_3072;
wire lut_f_3073;
wire lut_f_3074;
wire lut_f_3075;
wire lut_f_3076;
wire lut_f_3077;
wire lut_f_3078;
wire lut_f_3079;
wire lut_f_3080;
wire lut_f_3081;
wire lut_f_3082;
wire lut_f_3083;
wire lut_f_3084;
wire lut_f_3085;
wire lut_f_3086;
wire lut_f_3087;
wire lut_f_3088;
wire lut_f_3089;
wire lut_f_3090;
wire lut_f_3091;
wire lut_f_3092;
wire lut_f_3093;
wire lut_f_3094;
wire lut_f_3095;
wire lut_f_3096;
wire lut_f_3097;
wire lut_f_3098;
wire lut_f_3099;
wire lut_f_3100;
wire lut_f_3101;
wire lut_f_3102;
wire lut_f_3103;
wire lut_f_3104;
wire lut_f_3105;
wire lut_f_3106;
wire lut_f_3107;
wire lut_f_3108;
wire lut_f_3109;
wire lut_f_3110;
wire lut_f_3111;
wire lut_f_3112;
wire lut_f_3113;
wire lut_f_3114;
wire lut_f_3115;
wire lut_f_3116;
wire lut_f_3117;
wire lut_f_3118;
wire lut_f_3119;
wire lut_f_3120;
wire lut_f_3121;
wire lut_f_3122;
wire lut_f_3123;
wire lut_f_3124;
wire lut_f_3125;
wire lut_f_3126;
wire lut_f_3127;
wire lut_f_3128;
wire lut_f_3129;
wire lut_f_3130;
wire lut_f_3131;
wire lut_f_3132;
wire lut_f_3133;
wire lut_f_3134;
wire lut_f_3135;
wire lut_f_3136;
wire lut_f_3137;
wire lut_f_3138;
wire lut_f_3139;
wire lut_f_3140;
wire lut_f_3141;
wire lut_f_3142;
wire lut_f_3143;
wire lut_f_3144;
wire lut_f_3145;
wire lut_f_3146;
wire lut_f_3147;
wire lut_f_3148;
wire lut_f_3149;
wire lut_f_3150;
wire lut_f_3151;
wire lut_f_3152;
wire lut_f_3153;
wire lut_f_3154;
wire lut_f_3155;
wire lut_f_3156;
wire lut_f_3157;
wire lut_f_3158;
wire lut_f_3159;
wire lut_f_3160;
wire lut_f_3161;
wire lut_f_3162;
wire lut_f_3163;
wire lut_f_3164;
wire lut_f_3165;
wire lut_f_3166;
wire lut_f_3167;
wire lut_f_3168;
wire lut_f_3169;
wire lut_f_3170;
wire lut_f_3171;
wire lut_f_3172;
wire lut_f_3173;
wire lut_f_3174;
wire lut_f_3175;
wire lut_f_3176;
wire lut_f_3177;
wire lut_f_3178;
wire lut_f_3179;
wire lut_f_3180;
wire lut_f_3181;
wire lut_f_3182;
wire lut_f_3183;
wire lut_f_3184;
wire lut_f_3185;
wire lut_f_3186;
wire lut_f_3187;
wire lut_f_3188;
wire lut_f_3189;
wire lut_f_3190;
wire lut_f_3191;
wire lut_f_3192;
wire lut_f_3193;
wire lut_f_3194;
wire lut_f_3195;
wire lut_f_3196;
wire lut_f_3197;
wire lut_f_3198;
wire lut_f_3199;
wire [2:0] ram16s_inst_0_dout;
wire [2:0] ram16s_inst_1_dout;
wire [2:0] ram16s_inst_2_dout;
wire [2:0] ram16s_inst_3_dout;
wire [2:0] ram16s_inst_4_dout;
wire [2:0] ram16s_inst_5_dout;
wire [2:0] ram16s_inst_6_dout;
wire [2:0] ram16s_inst_7_dout;
wire [2:0] ram16s_inst_8_dout;
wire [2:0] ram16s_inst_9_dout;
wire [2:0] ram16s_inst_10_dout;
wire [2:0] ram16s_inst_11_dout;
wire [2:0] ram16s_inst_12_dout;
wire [2:0] ram16s_inst_13_dout;
wire [2:0] ram16s_inst_14_dout;
wire [2:0] ram16s_inst_15_dout;
wire [2:0] ram16s_inst_16_dout;
wire [2:0] ram16s_inst_17_dout;
wire [2:0] ram16s_inst_18_dout;
wire [2:0] ram16s_inst_19_dout;
wire [2:0] ram16s_inst_20_dout;
wire [2:0] ram16s_inst_21_dout;
wire [2:0] ram16s_inst_22_dout;
wire [2:0] ram16s_inst_23_dout;
wire [2:0] ram16s_inst_24_dout;
wire [2:0] ram16s_inst_25_dout;
wire [2:0] ram16s_inst_26_dout;
wire [2:0] ram16s_inst_27_dout;
wire [2:0] ram16s_inst_28_dout;
wire [2:0] ram16s_inst_29_dout;
wire [2:0] ram16s_inst_30_dout;
wire [2:0] ram16s_inst_31_dout;
wire [2:0] ram16s_inst_32_dout;
wire [2:0] ram16s_inst_33_dout;
wire [2:0] ram16s_inst_34_dout;
wire [2:0] ram16s_inst_35_dout;
wire [2:0] ram16s_inst_36_dout;
wire [2:0] ram16s_inst_37_dout;
wire [2:0] ram16s_inst_38_dout;
wire [2:0] ram16s_inst_39_dout;
wire [2:0] ram16s_inst_40_dout;
wire [2:0] ram16s_inst_41_dout;
wire [2:0] ram16s_inst_42_dout;
wire [2:0] ram16s_inst_43_dout;
wire [2:0] ram16s_inst_44_dout;
wire [2:0] ram16s_inst_45_dout;
wire [2:0] ram16s_inst_46_dout;
wire [2:0] ram16s_inst_47_dout;
wire [2:0] ram16s_inst_48_dout;
wire [2:0] ram16s_inst_49_dout;
wire [2:0] ram16s_inst_50_dout;
wire [2:0] ram16s_inst_51_dout;
wire [2:0] ram16s_inst_52_dout;
wire [2:0] ram16s_inst_53_dout;
wire [2:0] ram16s_inst_54_dout;
wire [2:0] ram16s_inst_55_dout;
wire [2:0] ram16s_inst_56_dout;
wire [2:0] ram16s_inst_57_dout;
wire [2:0] ram16s_inst_58_dout;
wire [2:0] ram16s_inst_59_dout;
wire [2:0] ram16s_inst_60_dout;
wire [2:0] ram16s_inst_61_dout;
wire [2:0] ram16s_inst_62_dout;
wire [2:0] ram16s_inst_63_dout;
wire [2:0] ram16s_inst_64_dout;
wire [2:0] ram16s_inst_65_dout;
wire [2:0] ram16s_inst_66_dout;
wire [2:0] ram16s_inst_67_dout;
wire [2:0] ram16s_inst_68_dout;
wire [2:0] ram16s_inst_69_dout;
wire [2:0] ram16s_inst_70_dout;
wire [2:0] ram16s_inst_71_dout;
wire [2:0] ram16s_inst_72_dout;
wire [2:0] ram16s_inst_73_dout;
wire [2:0] ram16s_inst_74_dout;
wire [2:0] ram16s_inst_75_dout;
wire [2:0] ram16s_inst_76_dout;
wire [2:0] ram16s_inst_77_dout;
wire [2:0] ram16s_inst_78_dout;
wire [2:0] ram16s_inst_79_dout;
wire [2:0] ram16s_inst_80_dout;
wire [2:0] ram16s_inst_81_dout;
wire [2:0] ram16s_inst_82_dout;
wire [2:0] ram16s_inst_83_dout;
wire [2:0] ram16s_inst_84_dout;
wire [2:0] ram16s_inst_85_dout;
wire [2:0] ram16s_inst_86_dout;
wire [2:0] ram16s_inst_87_dout;
wire [2:0] ram16s_inst_88_dout;
wire [2:0] ram16s_inst_89_dout;
wire [2:0] ram16s_inst_90_dout;
wire [2:0] ram16s_inst_91_dout;
wire [2:0] ram16s_inst_92_dout;
wire [2:0] ram16s_inst_93_dout;
wire [2:0] ram16s_inst_94_dout;
wire [2:0] ram16s_inst_95_dout;
wire [2:0] ram16s_inst_96_dout;
wire [2:0] ram16s_inst_97_dout;
wire [2:0] ram16s_inst_98_dout;
wire [2:0] ram16s_inst_99_dout;
wire [2:0] ram16s_inst_100_dout;
wire [2:0] ram16s_inst_101_dout;
wire [2:0] ram16s_inst_102_dout;
wire [2:0] ram16s_inst_103_dout;
wire [2:0] ram16s_inst_104_dout;
wire [2:0] ram16s_inst_105_dout;
wire [2:0] ram16s_inst_106_dout;
wire [2:0] ram16s_inst_107_dout;
wire [2:0] ram16s_inst_108_dout;
wire [2:0] ram16s_inst_109_dout;
wire [2:0] ram16s_inst_110_dout;
wire [2:0] ram16s_inst_111_dout;
wire [2:0] ram16s_inst_112_dout;
wire [2:0] ram16s_inst_113_dout;
wire [2:0] ram16s_inst_114_dout;
wire [2:0] ram16s_inst_115_dout;
wire [2:0] ram16s_inst_116_dout;
wire [2:0] ram16s_inst_117_dout;
wire [2:0] ram16s_inst_118_dout;
wire [2:0] ram16s_inst_119_dout;
wire [2:0] ram16s_inst_120_dout;
wire [2:0] ram16s_inst_121_dout;
wire [2:0] ram16s_inst_122_dout;
wire [2:0] ram16s_inst_123_dout;
wire [2:0] ram16s_inst_124_dout;
wire [2:0] ram16s_inst_125_dout;
wire [2:0] ram16s_inst_126_dout;
wire [2:0] ram16s_inst_127_dout;
wire [2:0] ram16s_inst_128_dout;
wire [2:0] ram16s_inst_129_dout;
wire [2:0] ram16s_inst_130_dout;
wire [2:0] ram16s_inst_131_dout;
wire [2:0] ram16s_inst_132_dout;
wire [2:0] ram16s_inst_133_dout;
wire [2:0] ram16s_inst_134_dout;
wire [2:0] ram16s_inst_135_dout;
wire [2:0] ram16s_inst_136_dout;
wire [2:0] ram16s_inst_137_dout;
wire [2:0] ram16s_inst_138_dout;
wire [2:0] ram16s_inst_139_dout;
wire [2:0] ram16s_inst_140_dout;
wire [2:0] ram16s_inst_141_dout;
wire [2:0] ram16s_inst_142_dout;
wire [2:0] ram16s_inst_143_dout;
wire [2:0] ram16s_inst_144_dout;
wire [2:0] ram16s_inst_145_dout;
wire [2:0] ram16s_inst_146_dout;
wire [2:0] ram16s_inst_147_dout;
wire [2:0] ram16s_inst_148_dout;
wire [2:0] ram16s_inst_149_dout;
wire [2:0] ram16s_inst_150_dout;
wire [2:0] ram16s_inst_151_dout;
wire [2:0] ram16s_inst_152_dout;
wire [2:0] ram16s_inst_153_dout;
wire [2:0] ram16s_inst_154_dout;
wire [2:0] ram16s_inst_155_dout;
wire [2:0] ram16s_inst_156_dout;
wire [2:0] ram16s_inst_157_dout;
wire [2:0] ram16s_inst_158_dout;
wire [2:0] ram16s_inst_159_dout;
wire [2:0] ram16s_inst_160_dout;
wire [2:0] ram16s_inst_161_dout;
wire [2:0] ram16s_inst_162_dout;
wire [2:0] ram16s_inst_163_dout;
wire [2:0] ram16s_inst_164_dout;
wire [2:0] ram16s_inst_165_dout;
wire [2:0] ram16s_inst_166_dout;
wire [2:0] ram16s_inst_167_dout;
wire [2:0] ram16s_inst_168_dout;
wire [2:0] ram16s_inst_169_dout;
wire [2:0] ram16s_inst_170_dout;
wire [2:0] ram16s_inst_171_dout;
wire [2:0] ram16s_inst_172_dout;
wire [2:0] ram16s_inst_173_dout;
wire [2:0] ram16s_inst_174_dout;
wire [2:0] ram16s_inst_175_dout;
wire [2:0] ram16s_inst_176_dout;
wire [2:0] ram16s_inst_177_dout;
wire [2:0] ram16s_inst_178_dout;
wire [2:0] ram16s_inst_179_dout;
wire [2:0] ram16s_inst_180_dout;
wire [2:0] ram16s_inst_181_dout;
wire [2:0] ram16s_inst_182_dout;
wire [2:0] ram16s_inst_183_dout;
wire [2:0] ram16s_inst_184_dout;
wire [2:0] ram16s_inst_185_dout;
wire [2:0] ram16s_inst_186_dout;
wire [2:0] ram16s_inst_187_dout;
wire [2:0] ram16s_inst_188_dout;
wire [2:0] ram16s_inst_189_dout;
wire [2:0] ram16s_inst_190_dout;
wire [2:0] ram16s_inst_191_dout;
wire [2:0] ram16s_inst_192_dout;
wire [2:0] ram16s_inst_193_dout;
wire [2:0] ram16s_inst_194_dout;
wire [2:0] ram16s_inst_195_dout;
wire [2:0] ram16s_inst_196_dout;
wire [2:0] ram16s_inst_197_dout;
wire [2:0] ram16s_inst_198_dout;
wire [2:0] ram16s_inst_199_dout;
wire [2:0] ram16s_inst_200_dout;
wire [2:0] ram16s_inst_201_dout;
wire [2:0] ram16s_inst_202_dout;
wire [2:0] ram16s_inst_203_dout;
wire [2:0] ram16s_inst_204_dout;
wire [2:0] ram16s_inst_205_dout;
wire [2:0] ram16s_inst_206_dout;
wire [2:0] ram16s_inst_207_dout;
wire [2:0] ram16s_inst_208_dout;
wire [2:0] ram16s_inst_209_dout;
wire [2:0] ram16s_inst_210_dout;
wire [2:0] ram16s_inst_211_dout;
wire [2:0] ram16s_inst_212_dout;
wire [2:0] ram16s_inst_213_dout;
wire [2:0] ram16s_inst_214_dout;
wire [2:0] ram16s_inst_215_dout;
wire [2:0] ram16s_inst_216_dout;
wire [2:0] ram16s_inst_217_dout;
wire [2:0] ram16s_inst_218_dout;
wire [2:0] ram16s_inst_219_dout;
wire [2:0] ram16s_inst_220_dout;
wire [2:0] ram16s_inst_221_dout;
wire [2:0] ram16s_inst_222_dout;
wire [2:0] ram16s_inst_223_dout;
wire [2:0] ram16s_inst_224_dout;
wire [2:0] ram16s_inst_225_dout;
wire [2:0] ram16s_inst_226_dout;
wire [2:0] ram16s_inst_227_dout;
wire [2:0] ram16s_inst_228_dout;
wire [2:0] ram16s_inst_229_dout;
wire [2:0] ram16s_inst_230_dout;
wire [2:0] ram16s_inst_231_dout;
wire [2:0] ram16s_inst_232_dout;
wire [2:0] ram16s_inst_233_dout;
wire [2:0] ram16s_inst_234_dout;
wire [2:0] ram16s_inst_235_dout;
wire [2:0] ram16s_inst_236_dout;
wire [2:0] ram16s_inst_237_dout;
wire [2:0] ram16s_inst_238_dout;
wire [2:0] ram16s_inst_239_dout;
wire [2:0] ram16s_inst_240_dout;
wire [2:0] ram16s_inst_241_dout;
wire [2:0] ram16s_inst_242_dout;
wire [2:0] ram16s_inst_243_dout;
wire [2:0] ram16s_inst_244_dout;
wire [2:0] ram16s_inst_245_dout;
wire [2:0] ram16s_inst_246_dout;
wire [2:0] ram16s_inst_247_dout;
wire [2:0] ram16s_inst_248_dout;
wire [2:0] ram16s_inst_249_dout;
wire [2:0] ram16s_inst_250_dout;
wire [2:0] ram16s_inst_251_dout;
wire [2:0] ram16s_inst_252_dout;
wire [2:0] ram16s_inst_253_dout;
wire [2:0] ram16s_inst_254_dout;
wire [2:0] ram16s_inst_255_dout;
wire [2:0] ram16s_inst_256_dout;
wire [2:0] ram16s_inst_257_dout;
wire [2:0] ram16s_inst_258_dout;
wire [2:0] ram16s_inst_259_dout;
wire [2:0] ram16s_inst_260_dout;
wire [2:0] ram16s_inst_261_dout;
wire [2:0] ram16s_inst_262_dout;
wire [2:0] ram16s_inst_263_dout;
wire [2:0] ram16s_inst_264_dout;
wire [2:0] ram16s_inst_265_dout;
wire [2:0] ram16s_inst_266_dout;
wire [2:0] ram16s_inst_267_dout;
wire [2:0] ram16s_inst_268_dout;
wire [2:0] ram16s_inst_269_dout;
wire [2:0] ram16s_inst_270_dout;
wire [2:0] ram16s_inst_271_dout;
wire [2:0] ram16s_inst_272_dout;
wire [2:0] ram16s_inst_273_dout;
wire [2:0] ram16s_inst_274_dout;
wire [2:0] ram16s_inst_275_dout;
wire [2:0] ram16s_inst_276_dout;
wire [2:0] ram16s_inst_277_dout;
wire [2:0] ram16s_inst_278_dout;
wire [2:0] ram16s_inst_279_dout;
wire [2:0] ram16s_inst_280_dout;
wire [2:0] ram16s_inst_281_dout;
wire [2:0] ram16s_inst_282_dout;
wire [2:0] ram16s_inst_283_dout;
wire [2:0] ram16s_inst_284_dout;
wire [2:0] ram16s_inst_285_dout;
wire [2:0] ram16s_inst_286_dout;
wire [2:0] ram16s_inst_287_dout;
wire [2:0] ram16s_inst_288_dout;
wire [2:0] ram16s_inst_289_dout;
wire [2:0] ram16s_inst_290_dout;
wire [2:0] ram16s_inst_291_dout;
wire [2:0] ram16s_inst_292_dout;
wire [2:0] ram16s_inst_293_dout;
wire [2:0] ram16s_inst_294_dout;
wire [2:0] ram16s_inst_295_dout;
wire [2:0] ram16s_inst_296_dout;
wire [2:0] ram16s_inst_297_dout;
wire [2:0] ram16s_inst_298_dout;
wire [2:0] ram16s_inst_299_dout;
wire [2:0] ram16s_inst_300_dout;
wire [2:0] ram16s_inst_301_dout;
wire [2:0] ram16s_inst_302_dout;
wire [2:0] ram16s_inst_303_dout;
wire [2:0] ram16s_inst_304_dout;
wire [2:0] ram16s_inst_305_dout;
wire [2:0] ram16s_inst_306_dout;
wire [2:0] ram16s_inst_307_dout;
wire [2:0] ram16s_inst_308_dout;
wire [2:0] ram16s_inst_309_dout;
wire [2:0] ram16s_inst_310_dout;
wire [2:0] ram16s_inst_311_dout;
wire [2:0] ram16s_inst_312_dout;
wire [2:0] ram16s_inst_313_dout;
wire [2:0] ram16s_inst_314_dout;
wire [2:0] ram16s_inst_315_dout;
wire [2:0] ram16s_inst_316_dout;
wire [2:0] ram16s_inst_317_dout;
wire [2:0] ram16s_inst_318_dout;
wire [2:0] ram16s_inst_319_dout;
wire [2:0] ram16s_inst_320_dout;
wire [2:0] ram16s_inst_321_dout;
wire [2:0] ram16s_inst_322_dout;
wire [2:0] ram16s_inst_323_dout;
wire [2:0] ram16s_inst_324_dout;
wire [2:0] ram16s_inst_325_dout;
wire [2:0] ram16s_inst_326_dout;
wire [2:0] ram16s_inst_327_dout;
wire [2:0] ram16s_inst_328_dout;
wire [2:0] ram16s_inst_329_dout;
wire [2:0] ram16s_inst_330_dout;
wire [2:0] ram16s_inst_331_dout;
wire [2:0] ram16s_inst_332_dout;
wire [2:0] ram16s_inst_333_dout;
wire [2:0] ram16s_inst_334_dout;
wire [2:0] ram16s_inst_335_dout;
wire [2:0] ram16s_inst_336_dout;
wire [2:0] ram16s_inst_337_dout;
wire [2:0] ram16s_inst_338_dout;
wire [2:0] ram16s_inst_339_dout;
wire [2:0] ram16s_inst_340_dout;
wire [2:0] ram16s_inst_341_dout;
wire [2:0] ram16s_inst_342_dout;
wire [2:0] ram16s_inst_343_dout;
wire [2:0] ram16s_inst_344_dout;
wire [2:0] ram16s_inst_345_dout;
wire [2:0] ram16s_inst_346_dout;
wire [2:0] ram16s_inst_347_dout;
wire [2:0] ram16s_inst_348_dout;
wire [2:0] ram16s_inst_349_dout;
wire [2:0] ram16s_inst_350_dout;
wire [2:0] ram16s_inst_351_dout;
wire [2:0] ram16s_inst_352_dout;
wire [2:0] ram16s_inst_353_dout;
wire [2:0] ram16s_inst_354_dout;
wire [2:0] ram16s_inst_355_dout;
wire [2:0] ram16s_inst_356_dout;
wire [2:0] ram16s_inst_357_dout;
wire [2:0] ram16s_inst_358_dout;
wire [2:0] ram16s_inst_359_dout;
wire [2:0] ram16s_inst_360_dout;
wire [2:0] ram16s_inst_361_dout;
wire [2:0] ram16s_inst_362_dout;
wire [2:0] ram16s_inst_363_dout;
wire [2:0] ram16s_inst_364_dout;
wire [2:0] ram16s_inst_365_dout;
wire [2:0] ram16s_inst_366_dout;
wire [2:0] ram16s_inst_367_dout;
wire [2:0] ram16s_inst_368_dout;
wire [2:0] ram16s_inst_369_dout;
wire [2:0] ram16s_inst_370_dout;
wire [2:0] ram16s_inst_371_dout;
wire [2:0] ram16s_inst_372_dout;
wire [2:0] ram16s_inst_373_dout;
wire [2:0] ram16s_inst_374_dout;
wire [2:0] ram16s_inst_375_dout;
wire [2:0] ram16s_inst_376_dout;
wire [2:0] ram16s_inst_377_dout;
wire [2:0] ram16s_inst_378_dout;
wire [2:0] ram16s_inst_379_dout;
wire [2:0] ram16s_inst_380_dout;
wire [2:0] ram16s_inst_381_dout;
wire [2:0] ram16s_inst_382_dout;
wire [2:0] ram16s_inst_383_dout;
wire [2:0] ram16s_inst_384_dout;
wire [2:0] ram16s_inst_385_dout;
wire [2:0] ram16s_inst_386_dout;
wire [2:0] ram16s_inst_387_dout;
wire [2:0] ram16s_inst_388_dout;
wire [2:0] ram16s_inst_389_dout;
wire [2:0] ram16s_inst_390_dout;
wire [2:0] ram16s_inst_391_dout;
wire [2:0] ram16s_inst_392_dout;
wire [2:0] ram16s_inst_393_dout;
wire [2:0] ram16s_inst_394_dout;
wire [2:0] ram16s_inst_395_dout;
wire [2:0] ram16s_inst_396_dout;
wire [2:0] ram16s_inst_397_dout;
wire [2:0] ram16s_inst_398_dout;
wire [2:0] ram16s_inst_399_dout;
wire [2:0] ram16s_inst_400_dout;
wire [2:0] ram16s_inst_401_dout;
wire [2:0] ram16s_inst_402_dout;
wire [2:0] ram16s_inst_403_dout;
wire [2:0] ram16s_inst_404_dout;
wire [2:0] ram16s_inst_405_dout;
wire [2:0] ram16s_inst_406_dout;
wire [2:0] ram16s_inst_407_dout;
wire [2:0] ram16s_inst_408_dout;
wire [2:0] ram16s_inst_409_dout;
wire [2:0] ram16s_inst_410_dout;
wire [2:0] ram16s_inst_411_dout;
wire [2:0] ram16s_inst_412_dout;
wire [2:0] ram16s_inst_413_dout;
wire [2:0] ram16s_inst_414_dout;
wire [2:0] ram16s_inst_415_dout;
wire [2:0] ram16s_inst_416_dout;
wire [2:0] ram16s_inst_417_dout;
wire [2:0] ram16s_inst_418_dout;
wire [2:0] ram16s_inst_419_dout;
wire [2:0] ram16s_inst_420_dout;
wire [2:0] ram16s_inst_421_dout;
wire [2:0] ram16s_inst_422_dout;
wire [2:0] ram16s_inst_423_dout;
wire [2:0] ram16s_inst_424_dout;
wire [2:0] ram16s_inst_425_dout;
wire [2:0] ram16s_inst_426_dout;
wire [2:0] ram16s_inst_427_dout;
wire [2:0] ram16s_inst_428_dout;
wire [2:0] ram16s_inst_429_dout;
wire [2:0] ram16s_inst_430_dout;
wire [2:0] ram16s_inst_431_dout;
wire [2:0] ram16s_inst_432_dout;
wire [2:0] ram16s_inst_433_dout;
wire [2:0] ram16s_inst_434_dout;
wire [2:0] ram16s_inst_435_dout;
wire [2:0] ram16s_inst_436_dout;
wire [2:0] ram16s_inst_437_dout;
wire [2:0] ram16s_inst_438_dout;
wire [2:0] ram16s_inst_439_dout;
wire [2:0] ram16s_inst_440_dout;
wire [2:0] ram16s_inst_441_dout;
wire [2:0] ram16s_inst_442_dout;
wire [2:0] ram16s_inst_443_dout;
wire [2:0] ram16s_inst_444_dout;
wire [2:0] ram16s_inst_445_dout;
wire [2:0] ram16s_inst_446_dout;
wire [2:0] ram16s_inst_447_dout;
wire [2:0] ram16s_inst_448_dout;
wire [2:0] ram16s_inst_449_dout;
wire [2:0] ram16s_inst_450_dout;
wire [2:0] ram16s_inst_451_dout;
wire [2:0] ram16s_inst_452_dout;
wire [2:0] ram16s_inst_453_dout;
wire [2:0] ram16s_inst_454_dout;
wire [2:0] ram16s_inst_455_dout;
wire [2:0] ram16s_inst_456_dout;
wire [2:0] ram16s_inst_457_dout;
wire [2:0] ram16s_inst_458_dout;
wire [2:0] ram16s_inst_459_dout;
wire [2:0] ram16s_inst_460_dout;
wire [2:0] ram16s_inst_461_dout;
wire [2:0] ram16s_inst_462_dout;
wire [2:0] ram16s_inst_463_dout;
wire [2:0] ram16s_inst_464_dout;
wire [2:0] ram16s_inst_465_dout;
wire [2:0] ram16s_inst_466_dout;
wire [2:0] ram16s_inst_467_dout;
wire [2:0] ram16s_inst_468_dout;
wire [2:0] ram16s_inst_469_dout;
wire [2:0] ram16s_inst_470_dout;
wire [2:0] ram16s_inst_471_dout;
wire [2:0] ram16s_inst_472_dout;
wire [2:0] ram16s_inst_473_dout;
wire [2:0] ram16s_inst_474_dout;
wire [2:0] ram16s_inst_475_dout;
wire [2:0] ram16s_inst_476_dout;
wire [2:0] ram16s_inst_477_dout;
wire [2:0] ram16s_inst_478_dout;
wire [2:0] ram16s_inst_479_dout;
wire [2:0] ram16s_inst_480_dout;
wire [2:0] ram16s_inst_481_dout;
wire [2:0] ram16s_inst_482_dout;
wire [2:0] ram16s_inst_483_dout;
wire [2:0] ram16s_inst_484_dout;
wire [2:0] ram16s_inst_485_dout;
wire [2:0] ram16s_inst_486_dout;
wire [2:0] ram16s_inst_487_dout;
wire [2:0] ram16s_inst_488_dout;
wire [2:0] ram16s_inst_489_dout;
wire [2:0] ram16s_inst_490_dout;
wire [2:0] ram16s_inst_491_dout;
wire [2:0] ram16s_inst_492_dout;
wire [2:0] ram16s_inst_493_dout;
wire [2:0] ram16s_inst_494_dout;
wire [2:0] ram16s_inst_495_dout;
wire [2:0] ram16s_inst_496_dout;
wire [2:0] ram16s_inst_497_dout;
wire [2:0] ram16s_inst_498_dout;
wire [2:0] ram16s_inst_499_dout;
wire [2:0] ram16s_inst_500_dout;
wire [2:0] ram16s_inst_501_dout;
wire [2:0] ram16s_inst_502_dout;
wire [2:0] ram16s_inst_503_dout;
wire [2:0] ram16s_inst_504_dout;
wire [2:0] ram16s_inst_505_dout;
wire [2:0] ram16s_inst_506_dout;
wire [2:0] ram16s_inst_507_dout;
wire [2:0] ram16s_inst_508_dout;
wire [2:0] ram16s_inst_509_dout;
wire [2:0] ram16s_inst_510_dout;
wire [2:0] ram16s_inst_511_dout;
wire [2:0] ram16s_inst_512_dout;
wire [2:0] ram16s_inst_513_dout;
wire [2:0] ram16s_inst_514_dout;
wire [2:0] ram16s_inst_515_dout;
wire [2:0] ram16s_inst_516_dout;
wire [2:0] ram16s_inst_517_dout;
wire [2:0] ram16s_inst_518_dout;
wire [2:0] ram16s_inst_519_dout;
wire [2:0] ram16s_inst_520_dout;
wire [2:0] ram16s_inst_521_dout;
wire [2:0] ram16s_inst_522_dout;
wire [2:0] ram16s_inst_523_dout;
wire [2:0] ram16s_inst_524_dout;
wire [2:0] ram16s_inst_525_dout;
wire [2:0] ram16s_inst_526_dout;
wire [2:0] ram16s_inst_527_dout;
wire [2:0] ram16s_inst_528_dout;
wire [2:0] ram16s_inst_529_dout;
wire [2:0] ram16s_inst_530_dout;
wire [2:0] ram16s_inst_531_dout;
wire [2:0] ram16s_inst_532_dout;
wire [2:0] ram16s_inst_533_dout;
wire [2:0] ram16s_inst_534_dout;
wire [2:0] ram16s_inst_535_dout;
wire [2:0] ram16s_inst_536_dout;
wire [2:0] ram16s_inst_537_dout;
wire [2:0] ram16s_inst_538_dout;
wire [2:0] ram16s_inst_539_dout;
wire [2:0] ram16s_inst_540_dout;
wire [2:0] ram16s_inst_541_dout;
wire [2:0] ram16s_inst_542_dout;
wire [2:0] ram16s_inst_543_dout;
wire [2:0] ram16s_inst_544_dout;
wire [2:0] ram16s_inst_545_dout;
wire [2:0] ram16s_inst_546_dout;
wire [2:0] ram16s_inst_547_dout;
wire [2:0] ram16s_inst_548_dout;
wire [2:0] ram16s_inst_549_dout;
wire [2:0] ram16s_inst_550_dout;
wire [2:0] ram16s_inst_551_dout;
wire [2:0] ram16s_inst_552_dout;
wire [2:0] ram16s_inst_553_dout;
wire [2:0] ram16s_inst_554_dout;
wire [2:0] ram16s_inst_555_dout;
wire [2:0] ram16s_inst_556_dout;
wire [2:0] ram16s_inst_557_dout;
wire [2:0] ram16s_inst_558_dout;
wire [2:0] ram16s_inst_559_dout;
wire [2:0] ram16s_inst_560_dout;
wire [2:0] ram16s_inst_561_dout;
wire [2:0] ram16s_inst_562_dout;
wire [2:0] ram16s_inst_563_dout;
wire [2:0] ram16s_inst_564_dout;
wire [2:0] ram16s_inst_565_dout;
wire [2:0] ram16s_inst_566_dout;
wire [2:0] ram16s_inst_567_dout;
wire [2:0] ram16s_inst_568_dout;
wire [2:0] ram16s_inst_569_dout;
wire [2:0] ram16s_inst_570_dout;
wire [2:0] ram16s_inst_571_dout;
wire [2:0] ram16s_inst_572_dout;
wire [2:0] ram16s_inst_573_dout;
wire [2:0] ram16s_inst_574_dout;
wire [2:0] ram16s_inst_575_dout;
wire [2:0] ram16s_inst_576_dout;
wire [2:0] ram16s_inst_577_dout;
wire [2:0] ram16s_inst_578_dout;
wire [2:0] ram16s_inst_579_dout;
wire [2:0] ram16s_inst_580_dout;
wire [2:0] ram16s_inst_581_dout;
wire [2:0] ram16s_inst_582_dout;
wire [2:0] ram16s_inst_583_dout;
wire [2:0] ram16s_inst_584_dout;
wire [2:0] ram16s_inst_585_dout;
wire [2:0] ram16s_inst_586_dout;
wire [2:0] ram16s_inst_587_dout;
wire [2:0] ram16s_inst_588_dout;
wire [2:0] ram16s_inst_589_dout;
wire [2:0] ram16s_inst_590_dout;
wire [2:0] ram16s_inst_591_dout;
wire [2:0] ram16s_inst_592_dout;
wire [2:0] ram16s_inst_593_dout;
wire [2:0] ram16s_inst_594_dout;
wire [2:0] ram16s_inst_595_dout;
wire [2:0] ram16s_inst_596_dout;
wire [2:0] ram16s_inst_597_dout;
wire [2:0] ram16s_inst_598_dout;
wire [2:0] ram16s_inst_599_dout;
wire [2:0] ram16s_inst_600_dout;
wire [2:0] ram16s_inst_601_dout;
wire [2:0] ram16s_inst_602_dout;
wire [2:0] ram16s_inst_603_dout;
wire [2:0] ram16s_inst_604_dout;
wire [2:0] ram16s_inst_605_dout;
wire [2:0] ram16s_inst_606_dout;
wire [2:0] ram16s_inst_607_dout;
wire [2:0] ram16s_inst_608_dout;
wire [2:0] ram16s_inst_609_dout;
wire [2:0] ram16s_inst_610_dout;
wire [2:0] ram16s_inst_611_dout;
wire [2:0] ram16s_inst_612_dout;
wire [2:0] ram16s_inst_613_dout;
wire [2:0] ram16s_inst_614_dout;
wire [2:0] ram16s_inst_615_dout;
wire [2:0] ram16s_inst_616_dout;
wire [2:0] ram16s_inst_617_dout;
wire [2:0] ram16s_inst_618_dout;
wire [2:0] ram16s_inst_619_dout;
wire [2:0] ram16s_inst_620_dout;
wire [2:0] ram16s_inst_621_dout;
wire [2:0] ram16s_inst_622_dout;
wire [2:0] ram16s_inst_623_dout;
wire [2:0] ram16s_inst_624_dout;
wire [2:0] ram16s_inst_625_dout;
wire [2:0] ram16s_inst_626_dout;
wire [2:0] ram16s_inst_627_dout;
wire [2:0] ram16s_inst_628_dout;
wire [2:0] ram16s_inst_629_dout;
wire [2:0] ram16s_inst_630_dout;
wire [2:0] ram16s_inst_631_dout;
wire [2:0] ram16s_inst_632_dout;
wire [2:0] ram16s_inst_633_dout;
wire [2:0] ram16s_inst_634_dout;
wire [2:0] ram16s_inst_635_dout;
wire [2:0] ram16s_inst_636_dout;
wire [2:0] ram16s_inst_637_dout;
wire [2:0] ram16s_inst_638_dout;
wire [2:0] ram16s_inst_639_dout;
wire [2:0] ram16s_inst_640_dout;
wire [2:0] ram16s_inst_641_dout;
wire [2:0] ram16s_inst_642_dout;
wire [2:0] ram16s_inst_643_dout;
wire [2:0] ram16s_inst_644_dout;
wire [2:0] ram16s_inst_645_dout;
wire [2:0] ram16s_inst_646_dout;
wire [2:0] ram16s_inst_647_dout;
wire [2:0] ram16s_inst_648_dout;
wire [2:0] ram16s_inst_649_dout;
wire [2:0] ram16s_inst_650_dout;
wire [2:0] ram16s_inst_651_dout;
wire [2:0] ram16s_inst_652_dout;
wire [2:0] ram16s_inst_653_dout;
wire [2:0] ram16s_inst_654_dout;
wire [2:0] ram16s_inst_655_dout;
wire [2:0] ram16s_inst_656_dout;
wire [2:0] ram16s_inst_657_dout;
wire [2:0] ram16s_inst_658_dout;
wire [2:0] ram16s_inst_659_dout;
wire [2:0] ram16s_inst_660_dout;
wire [2:0] ram16s_inst_661_dout;
wire [2:0] ram16s_inst_662_dout;
wire [2:0] ram16s_inst_663_dout;
wire [2:0] ram16s_inst_664_dout;
wire [2:0] ram16s_inst_665_dout;
wire [2:0] ram16s_inst_666_dout;
wire [2:0] ram16s_inst_667_dout;
wire [2:0] ram16s_inst_668_dout;
wire [2:0] ram16s_inst_669_dout;
wire [2:0] ram16s_inst_670_dout;
wire [2:0] ram16s_inst_671_dout;
wire [2:0] ram16s_inst_672_dout;
wire [2:0] ram16s_inst_673_dout;
wire [2:0] ram16s_inst_674_dout;
wire [2:0] ram16s_inst_675_dout;
wire [2:0] ram16s_inst_676_dout;
wire [2:0] ram16s_inst_677_dout;
wire [2:0] ram16s_inst_678_dout;
wire [2:0] ram16s_inst_679_dout;
wire [2:0] ram16s_inst_680_dout;
wire [2:0] ram16s_inst_681_dout;
wire [2:0] ram16s_inst_682_dout;
wire [2:0] ram16s_inst_683_dout;
wire [2:0] ram16s_inst_684_dout;
wire [2:0] ram16s_inst_685_dout;
wire [2:0] ram16s_inst_686_dout;
wire [2:0] ram16s_inst_687_dout;
wire [2:0] ram16s_inst_688_dout;
wire [2:0] ram16s_inst_689_dout;
wire [2:0] ram16s_inst_690_dout;
wire [2:0] ram16s_inst_691_dout;
wire [2:0] ram16s_inst_692_dout;
wire [2:0] ram16s_inst_693_dout;
wire [2:0] ram16s_inst_694_dout;
wire [2:0] ram16s_inst_695_dout;
wire [2:0] ram16s_inst_696_dout;
wire [2:0] ram16s_inst_697_dout;
wire [2:0] ram16s_inst_698_dout;
wire [2:0] ram16s_inst_699_dout;
wire [2:0] ram16s_inst_700_dout;
wire [2:0] ram16s_inst_701_dout;
wire [2:0] ram16s_inst_702_dout;
wire [2:0] ram16s_inst_703_dout;
wire [2:0] ram16s_inst_704_dout;
wire [2:0] ram16s_inst_705_dout;
wire [2:0] ram16s_inst_706_dout;
wire [2:0] ram16s_inst_707_dout;
wire [2:0] ram16s_inst_708_dout;
wire [2:0] ram16s_inst_709_dout;
wire [2:0] ram16s_inst_710_dout;
wire [2:0] ram16s_inst_711_dout;
wire [2:0] ram16s_inst_712_dout;
wire [2:0] ram16s_inst_713_dout;
wire [2:0] ram16s_inst_714_dout;
wire [2:0] ram16s_inst_715_dout;
wire [2:0] ram16s_inst_716_dout;
wire [2:0] ram16s_inst_717_dout;
wire [2:0] ram16s_inst_718_dout;
wire [2:0] ram16s_inst_719_dout;
wire [2:0] ram16s_inst_720_dout;
wire [2:0] ram16s_inst_721_dout;
wire [2:0] ram16s_inst_722_dout;
wire [2:0] ram16s_inst_723_dout;
wire [2:0] ram16s_inst_724_dout;
wire [2:0] ram16s_inst_725_dout;
wire [2:0] ram16s_inst_726_dout;
wire [2:0] ram16s_inst_727_dout;
wire [2:0] ram16s_inst_728_dout;
wire [2:0] ram16s_inst_729_dout;
wire [2:0] ram16s_inst_730_dout;
wire [2:0] ram16s_inst_731_dout;
wire [2:0] ram16s_inst_732_dout;
wire [2:0] ram16s_inst_733_dout;
wire [2:0] ram16s_inst_734_dout;
wire [2:0] ram16s_inst_735_dout;
wire [2:0] ram16s_inst_736_dout;
wire [2:0] ram16s_inst_737_dout;
wire [2:0] ram16s_inst_738_dout;
wire [2:0] ram16s_inst_739_dout;
wire [2:0] ram16s_inst_740_dout;
wire [2:0] ram16s_inst_741_dout;
wire [2:0] ram16s_inst_742_dout;
wire [2:0] ram16s_inst_743_dout;
wire [2:0] ram16s_inst_744_dout;
wire [2:0] ram16s_inst_745_dout;
wire [2:0] ram16s_inst_746_dout;
wire [2:0] ram16s_inst_747_dout;
wire [2:0] ram16s_inst_748_dout;
wire [2:0] ram16s_inst_749_dout;
wire [2:0] ram16s_inst_750_dout;
wire [2:0] ram16s_inst_751_dout;
wire [2:0] ram16s_inst_752_dout;
wire [2:0] ram16s_inst_753_dout;
wire [2:0] ram16s_inst_754_dout;
wire [2:0] ram16s_inst_755_dout;
wire [2:0] ram16s_inst_756_dout;
wire [2:0] ram16s_inst_757_dout;
wire [2:0] ram16s_inst_758_dout;
wire [2:0] ram16s_inst_759_dout;
wire [2:0] ram16s_inst_760_dout;
wire [2:0] ram16s_inst_761_dout;
wire [2:0] ram16s_inst_762_dout;
wire [2:0] ram16s_inst_763_dout;
wire [2:0] ram16s_inst_764_dout;
wire [2:0] ram16s_inst_765_dout;
wire [2:0] ram16s_inst_766_dout;
wire [2:0] ram16s_inst_767_dout;
wire [2:0] ram16s_inst_768_dout;
wire [2:0] ram16s_inst_769_dout;
wire [2:0] ram16s_inst_770_dout;
wire [2:0] ram16s_inst_771_dout;
wire [2:0] ram16s_inst_772_dout;
wire [2:0] ram16s_inst_773_dout;
wire [2:0] ram16s_inst_774_dout;
wire [2:0] ram16s_inst_775_dout;
wire [2:0] ram16s_inst_776_dout;
wire [2:0] ram16s_inst_777_dout;
wire [2:0] ram16s_inst_778_dout;
wire [2:0] ram16s_inst_779_dout;
wire [2:0] ram16s_inst_780_dout;
wire [2:0] ram16s_inst_781_dout;
wire [2:0] ram16s_inst_782_dout;
wire [2:0] ram16s_inst_783_dout;
wire [2:0] ram16s_inst_784_dout;
wire [2:0] ram16s_inst_785_dout;
wire [2:0] ram16s_inst_786_dout;
wire [2:0] ram16s_inst_787_dout;
wire [2:0] ram16s_inst_788_dout;
wire [2:0] ram16s_inst_789_dout;
wire [2:0] ram16s_inst_790_dout;
wire [2:0] ram16s_inst_791_dout;
wire [2:0] ram16s_inst_792_dout;
wire [2:0] ram16s_inst_793_dout;
wire [2:0] ram16s_inst_794_dout;
wire [2:0] ram16s_inst_795_dout;
wire [2:0] ram16s_inst_796_dout;
wire [2:0] ram16s_inst_797_dout;
wire [2:0] ram16s_inst_798_dout;
wire [2:0] ram16s_inst_799_dout;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_29;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_44;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_60;
wire mux_o_61;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_74;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_89;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_104;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_119;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_123;
wire mux_o_124;
wire mux_o_125;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_153;
wire mux_o_154;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_164;
wire mux_o_165;
wire mux_o_166;
wire mux_o_167;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_179;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_194;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_209;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_216;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_224;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_245;
wire mux_o_246;
wire mux_o_247;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_251;
wire mux_o_252;
wire mux_o_253;
wire mux_o_254;
wire mux_o_255;
wire mux_o_256;
wire mux_o_257;
wire mux_o_258;
wire mux_o_259;
wire mux_o_260;
wire mux_o_261;
wire mux_o_262;
wire mux_o_263;
wire mux_o_264;
wire mux_o_265;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_269;
wire mux_o_270;
wire mux_o_271;
wire mux_o_272;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_276;
wire mux_o_277;
wire mux_o_278;
wire mux_o_279;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_284;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_293;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_297;
wire mux_o_298;
wire mux_o_299;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_304;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_308;
wire mux_o_309;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_314;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_321;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_328;
wire mux_o_329;
wire mux_o_330;
wire mux_o_331;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_335;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_349;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_356;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_360;
wire mux_o_361;
wire mux_o_362;
wire mux_o_363;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_370;
wire mux_o_371;
wire mux_o_372;
wire mux_o_373;
wire mux_o_374;
wire mux_o_375;
wire mux_o_376;
wire mux_o_377;
wire mux_o_378;
wire mux_o_379;
wire mux_o_380;
wire mux_o_381;
wire mux_o_382;
wire mux_o_383;
wire mux_o_384;
wire mux_o_385;
wire mux_o_386;
wire mux_o_387;
wire mux_o_388;
wire mux_o_389;
wire mux_o_390;
wire mux_o_391;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_398;
wire mux_o_399;
wire mux_o_400;
wire mux_o_401;
wire mux_o_402;
wire mux_o_403;
wire mux_o_404;
wire mux_o_405;
wire mux_o_406;
wire mux_o_407;
wire mux_o_408;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_412;
wire mux_o_413;
wire mux_o_414;
wire mux_o_415;
wire mux_o_416;
wire mux_o_417;
wire mux_o_418;
wire mux_o_419;
wire mux_o_420;
wire mux_o_421;
wire mux_o_422;
wire mux_o_423;
wire mux_o_424;
wire mux_o_425;
wire mux_o_426;
wire mux_o_427;
wire mux_o_428;
wire mux_o_429;
wire mux_o_430;
wire mux_o_431;
wire mux_o_432;
wire mux_o_433;
wire mux_o_434;
wire mux_o_435;
wire mux_o_436;
wire mux_o_437;
wire mux_o_438;
wire mux_o_439;
wire mux_o_440;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire mux_o_447;
wire mux_o_448;
wire mux_o_449;
wire mux_o_450;
wire mux_o_451;
wire mux_o_452;
wire mux_o_453;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_459;
wire mux_o_460;
wire mux_o_461;
wire mux_o_462;
wire mux_o_463;
wire mux_o_464;
wire mux_o_465;
wire mux_o_466;
wire mux_o_467;
wire mux_o_468;
wire mux_o_469;
wire mux_o_470;
wire mux_o_471;
wire mux_o_472;
wire mux_o_473;
wire mux_o_474;
wire mux_o_475;
wire mux_o_476;
wire mux_o_477;
wire mux_o_478;
wire mux_o_479;
wire mux_o_480;
wire mux_o_481;
wire mux_o_482;
wire mux_o_483;
wire mux_o_484;
wire mux_o_485;
wire mux_o_486;
wire mux_o_487;
wire mux_o_488;
wire mux_o_489;
wire mux_o_490;
wire mux_o_491;
wire mux_o_492;
wire mux_o_493;
wire mux_o_494;
wire mux_o_495;
wire mux_o_496;
wire mux_o_497;
wire mux_o_498;
wire mux_o_499;
wire mux_o_500;
wire mux_o_501;
wire mux_o_502;
wire mux_o_503;
wire mux_o_504;
wire mux_o_505;
wire mux_o_506;
wire mux_o_507;
wire mux_o_508;
wire mux_o_509;
wire mux_o_510;
wire mux_o_511;
wire mux_o_512;
wire mux_o_513;
wire mux_o_514;
wire mux_o_515;
wire mux_o_516;
wire mux_o_517;
wire mux_o_518;
wire mux_o_519;
wire mux_o_520;
wire mux_o_521;
wire mux_o_522;
wire mux_o_523;
wire mux_o_524;
wire mux_o_525;
wire mux_o_526;
wire mux_o_527;
wire mux_o_528;
wire mux_o_529;
wire mux_o_530;
wire mux_o_531;
wire mux_o_532;
wire mux_o_533;
wire mux_o_534;
wire mux_o_535;
wire mux_o_536;
wire mux_o_537;
wire mux_o_538;
wire mux_o_539;
wire mux_o_540;
wire mux_o_541;
wire mux_o_542;
wire mux_o_543;
wire mux_o_544;
wire mux_o_545;
wire mux_o_546;
wire mux_o_547;
wire mux_o_548;
wire mux_o_549;
wire mux_o_550;
wire mux_o_551;
wire mux_o_552;
wire mux_o_553;
wire mux_o_554;
wire mux_o_555;
wire mux_o_556;
wire mux_o_557;
wire mux_o_558;
wire mux_o_559;
wire mux_o_560;
wire mux_o_561;
wire mux_o_562;
wire mux_o_563;
wire mux_o_564;
wire mux_o_565;
wire mux_o_566;
wire mux_o_567;
wire mux_o_568;
wire mux_o_569;
wire mux_o_570;
wire mux_o_571;
wire mux_o_572;
wire mux_o_573;
wire mux_o_574;
wire mux_o_575;
wire mux_o_576;
wire mux_o_577;
wire mux_o_578;
wire mux_o_579;
wire mux_o_580;
wire mux_o_581;
wire mux_o_582;
wire mux_o_583;
wire mux_o_584;
wire mux_o_585;
wire mux_o_586;
wire mux_o_587;
wire mux_o_588;
wire mux_o_589;
wire mux_o_590;
wire mux_o_591;
wire mux_o_592;
wire mux_o_593;
wire mux_o_594;
wire mux_o_595;
wire mux_o_596;
wire mux_o_597;
wire mux_o_598;
wire mux_o_599;
wire mux_o_600;
wire mux_o_601;
wire mux_o_602;
wire mux_o_603;
wire mux_o_604;
wire mux_o_605;
wire mux_o_606;
wire mux_o_607;
wire mux_o_608;
wire mux_o_609;
wire mux_o_610;
wire mux_o_611;
wire mux_o_612;
wire mux_o_613;
wire mux_o_614;
wire mux_o_615;
wire mux_o_616;
wire mux_o_617;
wire mux_o_618;
wire mux_o_619;
wire mux_o_620;
wire mux_o_621;
wire mux_o_622;
wire mux_o_623;
wire mux_o_624;
wire mux_o_625;
wire mux_o_626;
wire mux_o_627;
wire mux_o_628;
wire mux_o_629;
wire mux_o_630;
wire mux_o_631;
wire mux_o_632;
wire mux_o_633;
wire mux_o_634;
wire mux_o_635;
wire mux_o_636;
wire mux_o_637;
wire mux_o_638;
wire mux_o_639;
wire mux_o_640;
wire mux_o_641;
wire mux_o_642;
wire mux_o_643;
wire mux_o_644;
wire mux_o_645;
wire mux_o_646;
wire mux_o_647;
wire mux_o_648;
wire mux_o_649;
wire mux_o_650;
wire mux_o_651;
wire mux_o_652;
wire mux_o_653;
wire mux_o_654;
wire mux_o_655;
wire mux_o_656;
wire mux_o_657;
wire mux_o_658;
wire mux_o_659;
wire mux_o_660;
wire mux_o_661;
wire mux_o_662;
wire mux_o_663;
wire mux_o_664;
wire mux_o_665;
wire mux_o_666;
wire mux_o_667;
wire mux_o_668;
wire mux_o_669;
wire mux_o_670;
wire mux_o_671;
wire mux_o_672;
wire mux_o_673;
wire mux_o_674;
wire mux_o_675;
wire mux_o_676;
wire mux_o_677;
wire mux_o_678;
wire mux_o_679;
wire mux_o_680;
wire mux_o_681;
wire mux_o_682;
wire mux_o_683;
wire mux_o_684;
wire mux_o_685;
wire mux_o_686;
wire mux_o_687;
wire mux_o_688;
wire mux_o_689;
wire mux_o_690;
wire mux_o_691;
wire mux_o_692;
wire mux_o_693;
wire mux_o_694;
wire mux_o_695;
wire mux_o_696;
wire mux_o_697;
wire mux_o_698;
wire mux_o_699;
wire mux_o_700;
wire mux_o_701;
wire mux_o_702;
wire mux_o_703;
wire mux_o_704;
wire mux_o_705;
wire mux_o_706;
wire mux_o_707;
wire mux_o_708;
wire mux_o_709;
wire mux_o_710;
wire mux_o_711;
wire mux_o_712;
wire mux_o_713;
wire mux_o_714;
wire mux_o_715;
wire mux_o_716;
wire mux_o_717;
wire mux_o_718;
wire mux_o_719;
wire mux_o_720;
wire mux_o_721;
wire mux_o_722;
wire mux_o_723;
wire mux_o_724;
wire mux_o_725;
wire mux_o_726;
wire mux_o_727;
wire mux_o_728;
wire mux_o_729;
wire mux_o_730;
wire mux_o_731;
wire mux_o_732;
wire mux_o_733;
wire mux_o_734;
wire mux_o_735;
wire mux_o_736;
wire mux_o_737;
wire mux_o_738;
wire mux_o_739;
wire mux_o_740;
wire mux_o_741;
wire mux_o_742;
wire mux_o_743;
wire mux_o_744;
wire mux_o_745;
wire mux_o_746;
wire mux_o_747;
wire mux_o_748;
wire mux_o_749;
wire mux_o_750;
wire mux_o_751;
wire mux_o_752;
wire mux_o_753;
wire mux_o_754;
wire mux_o_755;
wire mux_o_756;
wire mux_o_757;
wire mux_o_758;
wire mux_o_759;
wire mux_o_760;
wire mux_o_761;
wire mux_o_762;
wire mux_o_763;
wire mux_o_764;
wire mux_o_765;
wire mux_o_766;
wire mux_o_767;
wire mux_o_768;
wire mux_o_769;
wire mux_o_770;
wire mux_o_771;
wire mux_o_772;
wire mux_o_773;
wire mux_o_774;
wire mux_o_775;
wire mux_o_776;
wire mux_o_777;
wire mux_o_778;
wire mux_o_779;
wire mux_o_780;
wire mux_o_781;
wire mux_o_782;
wire mux_o_783;
wire mux_o_784;
wire mux_o_785;
wire mux_o_786;
wire mux_o_788;
wire mux_o_789;
wire mux_o_790;
wire mux_o_791;
wire mux_o_792;
wire mux_o_793;
wire mux_o_795;
wire mux_o_796;
wire mux_o_797;
wire mux_o_799;
wire mux_o_800;
wire mux_o_802;
wire mux_o_803;
wire mux_o_804;
wire mux_o_805;
wire mux_o_806;
wire mux_o_807;
wire mux_o_808;
wire mux_o_809;
wire mux_o_810;
wire mux_o_811;
wire mux_o_812;
wire mux_o_813;
wire mux_o_814;
wire mux_o_815;
wire mux_o_816;
wire mux_o_817;
wire mux_o_818;
wire mux_o_819;
wire mux_o_820;
wire mux_o_821;
wire mux_o_822;
wire mux_o_823;
wire mux_o_824;
wire mux_o_825;
wire mux_o_826;
wire mux_o_827;
wire mux_o_828;
wire mux_o_829;
wire mux_o_830;
wire mux_o_831;
wire mux_o_832;
wire mux_o_833;
wire mux_o_834;
wire mux_o_835;
wire mux_o_836;
wire mux_o_837;
wire mux_o_838;
wire mux_o_839;
wire mux_o_840;
wire mux_o_841;
wire mux_o_842;
wire mux_o_843;
wire mux_o_844;
wire mux_o_845;
wire mux_o_846;
wire mux_o_847;
wire mux_o_848;
wire mux_o_849;
wire mux_o_850;
wire mux_o_851;
wire mux_o_852;
wire mux_o_853;
wire mux_o_854;
wire mux_o_855;
wire mux_o_856;
wire mux_o_857;
wire mux_o_858;
wire mux_o_859;
wire mux_o_860;
wire mux_o_861;
wire mux_o_862;
wire mux_o_863;
wire mux_o_864;
wire mux_o_865;
wire mux_o_866;
wire mux_o_867;
wire mux_o_868;
wire mux_o_869;
wire mux_o_870;
wire mux_o_871;
wire mux_o_872;
wire mux_o_873;
wire mux_o_874;
wire mux_o_875;
wire mux_o_876;
wire mux_o_877;
wire mux_o_878;
wire mux_o_879;
wire mux_o_880;
wire mux_o_881;
wire mux_o_882;
wire mux_o_883;
wire mux_o_884;
wire mux_o_885;
wire mux_o_886;
wire mux_o_887;
wire mux_o_888;
wire mux_o_889;
wire mux_o_890;
wire mux_o_891;
wire mux_o_892;
wire mux_o_893;
wire mux_o_894;
wire mux_o_895;
wire mux_o_896;
wire mux_o_897;
wire mux_o_898;
wire mux_o_899;
wire mux_o_900;
wire mux_o_901;
wire mux_o_902;
wire mux_o_903;
wire mux_o_904;
wire mux_o_905;
wire mux_o_906;
wire mux_o_907;
wire mux_o_908;
wire mux_o_909;
wire mux_o_910;
wire mux_o_911;
wire mux_o_912;
wire mux_o_913;
wire mux_o_914;
wire mux_o_915;
wire mux_o_916;
wire mux_o_917;
wire mux_o_918;
wire mux_o_919;
wire mux_o_920;
wire mux_o_921;
wire mux_o_922;
wire mux_o_923;
wire mux_o_924;
wire mux_o_925;
wire mux_o_926;
wire mux_o_927;
wire mux_o_928;
wire mux_o_929;
wire mux_o_930;
wire mux_o_931;
wire mux_o_932;
wire mux_o_933;
wire mux_o_934;
wire mux_o_935;
wire mux_o_936;
wire mux_o_937;
wire mux_o_938;
wire mux_o_939;
wire mux_o_940;
wire mux_o_941;
wire mux_o_942;
wire mux_o_943;
wire mux_o_944;
wire mux_o_945;
wire mux_o_946;
wire mux_o_947;
wire mux_o_948;
wire mux_o_949;
wire mux_o_950;
wire mux_o_951;
wire mux_o_952;
wire mux_o_953;
wire mux_o_954;
wire mux_o_955;
wire mux_o_956;
wire mux_o_957;
wire mux_o_958;
wire mux_o_959;
wire mux_o_960;
wire mux_o_961;
wire mux_o_962;
wire mux_o_963;
wire mux_o_964;
wire mux_o_965;
wire mux_o_966;
wire mux_o_967;
wire mux_o_968;
wire mux_o_969;
wire mux_o_970;
wire mux_o_971;
wire mux_o_972;
wire mux_o_973;
wire mux_o_974;
wire mux_o_975;
wire mux_o_976;
wire mux_o_977;
wire mux_o_978;
wire mux_o_979;
wire mux_o_980;
wire mux_o_981;
wire mux_o_982;
wire mux_o_983;
wire mux_o_984;
wire mux_o_985;
wire mux_o_986;
wire mux_o_987;
wire mux_o_988;
wire mux_o_989;
wire mux_o_990;
wire mux_o_991;
wire mux_o_992;
wire mux_o_993;
wire mux_o_994;
wire mux_o_995;
wire mux_o_996;
wire mux_o_997;
wire mux_o_998;
wire mux_o_999;
wire mux_o_1000;
wire mux_o_1001;
wire mux_o_1002;
wire mux_o_1003;
wire mux_o_1004;
wire mux_o_1005;
wire mux_o_1006;
wire mux_o_1007;
wire mux_o_1008;
wire mux_o_1009;
wire mux_o_1010;
wire mux_o_1011;
wire mux_o_1012;
wire mux_o_1013;
wire mux_o_1014;
wire mux_o_1015;
wire mux_o_1016;
wire mux_o_1017;
wire mux_o_1018;
wire mux_o_1019;
wire mux_o_1020;
wire mux_o_1021;
wire mux_o_1022;
wire mux_o_1023;
wire mux_o_1024;
wire mux_o_1025;
wire mux_o_1026;
wire mux_o_1027;
wire mux_o_1028;
wire mux_o_1029;
wire mux_o_1030;
wire mux_o_1031;
wire mux_o_1032;
wire mux_o_1033;
wire mux_o_1034;
wire mux_o_1035;
wire mux_o_1036;
wire mux_o_1037;
wire mux_o_1038;
wire mux_o_1039;
wire mux_o_1040;
wire mux_o_1041;
wire mux_o_1042;
wire mux_o_1043;
wire mux_o_1044;
wire mux_o_1045;
wire mux_o_1046;
wire mux_o_1047;
wire mux_o_1048;
wire mux_o_1049;
wire mux_o_1050;
wire mux_o_1051;
wire mux_o_1052;
wire mux_o_1053;
wire mux_o_1054;
wire mux_o_1055;
wire mux_o_1056;
wire mux_o_1057;
wire mux_o_1058;
wire mux_o_1059;
wire mux_o_1060;
wire mux_o_1061;
wire mux_o_1062;
wire mux_o_1063;
wire mux_o_1064;
wire mux_o_1065;
wire mux_o_1066;
wire mux_o_1067;
wire mux_o_1068;
wire mux_o_1069;
wire mux_o_1070;
wire mux_o_1071;
wire mux_o_1072;
wire mux_o_1073;
wire mux_o_1074;
wire mux_o_1075;
wire mux_o_1076;
wire mux_o_1077;
wire mux_o_1078;
wire mux_o_1079;
wire mux_o_1080;
wire mux_o_1081;
wire mux_o_1082;
wire mux_o_1083;
wire mux_o_1084;
wire mux_o_1085;
wire mux_o_1086;
wire mux_o_1087;
wire mux_o_1088;
wire mux_o_1089;
wire mux_o_1090;
wire mux_o_1091;
wire mux_o_1092;
wire mux_o_1093;
wire mux_o_1094;
wire mux_o_1095;
wire mux_o_1096;
wire mux_o_1097;
wire mux_o_1098;
wire mux_o_1099;
wire mux_o_1100;
wire mux_o_1101;
wire mux_o_1102;
wire mux_o_1103;
wire mux_o_1104;
wire mux_o_1105;
wire mux_o_1106;
wire mux_o_1107;
wire mux_o_1108;
wire mux_o_1109;
wire mux_o_1110;
wire mux_o_1111;
wire mux_o_1112;
wire mux_o_1113;
wire mux_o_1114;
wire mux_o_1115;
wire mux_o_1116;
wire mux_o_1117;
wire mux_o_1118;
wire mux_o_1119;
wire mux_o_1120;
wire mux_o_1121;
wire mux_o_1122;
wire mux_o_1123;
wire mux_o_1124;
wire mux_o_1125;
wire mux_o_1126;
wire mux_o_1127;
wire mux_o_1128;
wire mux_o_1129;
wire mux_o_1130;
wire mux_o_1131;
wire mux_o_1132;
wire mux_o_1133;
wire mux_o_1134;
wire mux_o_1135;
wire mux_o_1136;
wire mux_o_1137;
wire mux_o_1138;
wire mux_o_1139;
wire mux_o_1140;
wire mux_o_1141;
wire mux_o_1142;
wire mux_o_1143;
wire mux_o_1144;
wire mux_o_1145;
wire mux_o_1146;
wire mux_o_1147;
wire mux_o_1148;
wire mux_o_1149;
wire mux_o_1150;
wire mux_o_1151;
wire mux_o_1152;
wire mux_o_1153;
wire mux_o_1154;
wire mux_o_1155;
wire mux_o_1156;
wire mux_o_1157;
wire mux_o_1158;
wire mux_o_1159;
wire mux_o_1160;
wire mux_o_1161;
wire mux_o_1162;
wire mux_o_1163;
wire mux_o_1164;
wire mux_o_1165;
wire mux_o_1166;
wire mux_o_1167;
wire mux_o_1168;
wire mux_o_1169;
wire mux_o_1170;
wire mux_o_1171;
wire mux_o_1172;
wire mux_o_1173;
wire mux_o_1174;
wire mux_o_1175;
wire mux_o_1176;
wire mux_o_1177;
wire mux_o_1178;
wire mux_o_1179;
wire mux_o_1180;
wire mux_o_1181;
wire mux_o_1182;
wire mux_o_1183;
wire mux_o_1184;
wire mux_o_1185;
wire mux_o_1186;
wire mux_o_1187;
wire mux_o_1188;
wire mux_o_1189;
wire mux_o_1190;
wire mux_o_1191;
wire mux_o_1192;
wire mux_o_1193;
wire mux_o_1194;
wire mux_o_1195;
wire mux_o_1196;
wire mux_o_1197;
wire mux_o_1198;
wire mux_o_1199;
wire mux_o_1200;
wire mux_o_1201;
wire mux_o_1202;
wire mux_o_1203;
wire mux_o_1204;
wire mux_o_1205;
wire mux_o_1206;
wire mux_o_1207;
wire mux_o_1208;
wire mux_o_1209;
wire mux_o_1210;
wire mux_o_1211;
wire mux_o_1212;
wire mux_o_1213;
wire mux_o_1214;
wire mux_o_1215;
wire mux_o_1216;
wire mux_o_1217;
wire mux_o_1218;
wire mux_o_1219;
wire mux_o_1220;
wire mux_o_1221;
wire mux_o_1222;
wire mux_o_1223;
wire mux_o_1224;
wire mux_o_1225;
wire mux_o_1226;
wire mux_o_1227;
wire mux_o_1228;
wire mux_o_1229;
wire mux_o_1230;
wire mux_o_1231;
wire mux_o_1232;
wire mux_o_1233;
wire mux_o_1234;
wire mux_o_1235;
wire mux_o_1236;
wire mux_o_1237;
wire mux_o_1238;
wire mux_o_1239;
wire mux_o_1240;
wire mux_o_1241;
wire mux_o_1242;
wire mux_o_1243;
wire mux_o_1244;
wire mux_o_1245;
wire mux_o_1246;
wire mux_o_1247;
wire mux_o_1248;
wire mux_o_1249;
wire mux_o_1250;
wire mux_o_1251;
wire mux_o_1252;
wire mux_o_1253;
wire mux_o_1254;
wire mux_o_1255;
wire mux_o_1256;
wire mux_o_1257;
wire mux_o_1258;
wire mux_o_1259;
wire mux_o_1260;
wire mux_o_1261;
wire mux_o_1262;
wire mux_o_1263;
wire mux_o_1264;
wire mux_o_1265;
wire mux_o_1266;
wire mux_o_1267;
wire mux_o_1268;
wire mux_o_1269;
wire mux_o_1270;
wire mux_o_1271;
wire mux_o_1272;
wire mux_o_1273;
wire mux_o_1274;
wire mux_o_1275;
wire mux_o_1276;
wire mux_o_1277;
wire mux_o_1278;
wire mux_o_1279;
wire mux_o_1280;
wire mux_o_1281;
wire mux_o_1282;
wire mux_o_1283;
wire mux_o_1284;
wire mux_o_1285;
wire mux_o_1286;
wire mux_o_1287;
wire mux_o_1288;
wire mux_o_1289;
wire mux_o_1290;
wire mux_o_1291;
wire mux_o_1292;
wire mux_o_1293;
wire mux_o_1294;
wire mux_o_1295;
wire mux_o_1296;
wire mux_o_1297;
wire mux_o_1298;
wire mux_o_1299;
wire mux_o_1300;
wire mux_o_1301;
wire mux_o_1302;
wire mux_o_1303;
wire mux_o_1304;
wire mux_o_1305;
wire mux_o_1306;
wire mux_o_1307;
wire mux_o_1308;
wire mux_o_1309;
wire mux_o_1310;
wire mux_o_1311;
wire mux_o_1312;
wire mux_o_1313;
wire mux_o_1314;
wire mux_o_1315;
wire mux_o_1316;
wire mux_o_1317;
wire mux_o_1318;
wire mux_o_1319;
wire mux_o_1320;
wire mux_o_1321;
wire mux_o_1322;
wire mux_o_1323;
wire mux_o_1324;
wire mux_o_1325;
wire mux_o_1326;
wire mux_o_1327;
wire mux_o_1328;
wire mux_o_1329;
wire mux_o_1330;
wire mux_o_1331;
wire mux_o_1332;
wire mux_o_1333;
wire mux_o_1334;
wire mux_o_1335;
wire mux_o_1336;
wire mux_o_1337;
wire mux_o_1338;
wire mux_o_1339;
wire mux_o_1340;
wire mux_o_1341;
wire mux_o_1342;
wire mux_o_1343;
wire mux_o_1344;
wire mux_o_1345;
wire mux_o_1346;
wire mux_o_1347;
wire mux_o_1348;
wire mux_o_1349;
wire mux_o_1350;
wire mux_o_1351;
wire mux_o_1352;
wire mux_o_1353;
wire mux_o_1354;
wire mux_o_1355;
wire mux_o_1356;
wire mux_o_1357;
wire mux_o_1358;
wire mux_o_1359;
wire mux_o_1360;
wire mux_o_1361;
wire mux_o_1362;
wire mux_o_1363;
wire mux_o_1364;
wire mux_o_1365;
wire mux_o_1366;
wire mux_o_1367;
wire mux_o_1368;
wire mux_o_1369;
wire mux_o_1370;
wire mux_o_1371;
wire mux_o_1372;
wire mux_o_1373;
wire mux_o_1374;
wire mux_o_1375;
wire mux_o_1376;
wire mux_o_1377;
wire mux_o_1378;
wire mux_o_1379;
wire mux_o_1380;
wire mux_o_1381;
wire mux_o_1382;
wire mux_o_1383;
wire mux_o_1384;
wire mux_o_1385;
wire mux_o_1386;
wire mux_o_1387;
wire mux_o_1388;
wire mux_o_1389;
wire mux_o_1390;
wire mux_o_1391;
wire mux_o_1392;
wire mux_o_1393;
wire mux_o_1394;
wire mux_o_1395;
wire mux_o_1396;
wire mux_o_1397;
wire mux_o_1398;
wire mux_o_1399;
wire mux_o_1400;
wire mux_o_1401;
wire mux_o_1402;
wire mux_o_1403;
wire mux_o_1404;
wire mux_o_1405;
wire mux_o_1406;
wire mux_o_1407;
wire mux_o_1408;
wire mux_o_1409;
wire mux_o_1410;
wire mux_o_1411;
wire mux_o_1412;
wire mux_o_1413;
wire mux_o_1414;
wire mux_o_1415;
wire mux_o_1416;
wire mux_o_1417;
wire mux_o_1418;
wire mux_o_1419;
wire mux_o_1420;
wire mux_o_1421;
wire mux_o_1422;
wire mux_o_1423;
wire mux_o_1424;
wire mux_o_1425;
wire mux_o_1426;
wire mux_o_1427;
wire mux_o_1428;
wire mux_o_1429;
wire mux_o_1430;
wire mux_o_1431;
wire mux_o_1432;
wire mux_o_1433;
wire mux_o_1434;
wire mux_o_1435;
wire mux_o_1436;
wire mux_o_1437;
wire mux_o_1438;
wire mux_o_1439;
wire mux_o_1440;
wire mux_o_1441;
wire mux_o_1442;
wire mux_o_1443;
wire mux_o_1444;
wire mux_o_1445;
wire mux_o_1446;
wire mux_o_1447;
wire mux_o_1448;
wire mux_o_1449;
wire mux_o_1450;
wire mux_o_1451;
wire mux_o_1452;
wire mux_o_1453;
wire mux_o_1454;
wire mux_o_1455;
wire mux_o_1456;
wire mux_o_1457;
wire mux_o_1458;
wire mux_o_1459;
wire mux_o_1460;
wire mux_o_1461;
wire mux_o_1462;
wire mux_o_1463;
wire mux_o_1464;
wire mux_o_1465;
wire mux_o_1466;
wire mux_o_1467;
wire mux_o_1468;
wire mux_o_1469;
wire mux_o_1470;
wire mux_o_1471;
wire mux_o_1472;
wire mux_o_1473;
wire mux_o_1474;
wire mux_o_1475;
wire mux_o_1476;
wire mux_o_1477;
wire mux_o_1478;
wire mux_o_1479;
wire mux_o_1480;
wire mux_o_1481;
wire mux_o_1482;
wire mux_o_1483;
wire mux_o_1484;
wire mux_o_1485;
wire mux_o_1486;
wire mux_o_1487;
wire mux_o_1488;
wire mux_o_1489;
wire mux_o_1490;
wire mux_o_1491;
wire mux_o_1492;
wire mux_o_1493;
wire mux_o_1494;
wire mux_o_1495;
wire mux_o_1496;
wire mux_o_1497;
wire mux_o_1498;
wire mux_o_1499;
wire mux_o_1500;
wire mux_o_1501;
wire mux_o_1502;
wire mux_o_1503;
wire mux_o_1504;
wire mux_o_1505;
wire mux_o_1506;
wire mux_o_1507;
wire mux_o_1508;
wire mux_o_1509;
wire mux_o_1510;
wire mux_o_1511;
wire mux_o_1512;
wire mux_o_1513;
wire mux_o_1514;
wire mux_o_1515;
wire mux_o_1516;
wire mux_o_1517;
wire mux_o_1518;
wire mux_o_1519;
wire mux_o_1520;
wire mux_o_1521;
wire mux_o_1522;
wire mux_o_1523;
wire mux_o_1524;
wire mux_o_1525;
wire mux_o_1526;
wire mux_o_1527;
wire mux_o_1528;
wire mux_o_1529;
wire mux_o_1530;
wire mux_o_1531;
wire mux_o_1532;
wire mux_o_1533;
wire mux_o_1534;
wire mux_o_1535;
wire mux_o_1536;
wire mux_o_1537;
wire mux_o_1538;
wire mux_o_1539;
wire mux_o_1540;
wire mux_o_1541;
wire mux_o_1542;
wire mux_o_1543;
wire mux_o_1544;
wire mux_o_1545;
wire mux_o_1546;
wire mux_o_1547;
wire mux_o_1548;
wire mux_o_1549;
wire mux_o_1550;
wire mux_o_1551;
wire mux_o_1552;
wire mux_o_1553;
wire mux_o_1554;
wire mux_o_1555;
wire mux_o_1556;
wire mux_o_1557;
wire mux_o_1558;
wire mux_o_1559;
wire mux_o_1560;
wire mux_o_1561;
wire mux_o_1562;
wire mux_o_1563;
wire mux_o_1564;
wire mux_o_1565;
wire mux_o_1566;
wire mux_o_1567;
wire mux_o_1568;
wire mux_o_1569;
wire mux_o_1570;
wire mux_o_1571;
wire mux_o_1572;
wire mux_o_1573;
wire mux_o_1574;
wire mux_o_1575;
wire mux_o_1576;
wire mux_o_1577;
wire mux_o_1578;
wire mux_o_1579;
wire mux_o_1580;
wire mux_o_1581;
wire mux_o_1582;
wire mux_o_1583;
wire mux_o_1584;
wire mux_o_1585;
wire mux_o_1586;
wire mux_o_1587;
wire mux_o_1588;
wire mux_o_1590;
wire mux_o_1591;
wire mux_o_1592;
wire mux_o_1593;
wire mux_o_1594;
wire mux_o_1595;
wire mux_o_1597;
wire mux_o_1598;
wire mux_o_1599;
wire mux_o_1601;
wire mux_o_1602;
wire mux_o_1604;
wire mux_o_1605;
wire mux_o_1606;
wire mux_o_1607;
wire mux_o_1608;
wire mux_o_1609;
wire mux_o_1610;
wire mux_o_1611;
wire mux_o_1612;
wire mux_o_1613;
wire mux_o_1614;
wire mux_o_1615;
wire mux_o_1616;
wire mux_o_1617;
wire mux_o_1618;
wire mux_o_1619;
wire mux_o_1620;
wire mux_o_1621;
wire mux_o_1622;
wire mux_o_1623;
wire mux_o_1624;
wire mux_o_1625;
wire mux_o_1626;
wire mux_o_1627;
wire mux_o_1628;
wire mux_o_1629;
wire mux_o_1630;
wire mux_o_1631;
wire mux_o_1632;
wire mux_o_1633;
wire mux_o_1634;
wire mux_o_1635;
wire mux_o_1636;
wire mux_o_1637;
wire mux_o_1638;
wire mux_o_1639;
wire mux_o_1640;
wire mux_o_1641;
wire mux_o_1642;
wire mux_o_1643;
wire mux_o_1644;
wire mux_o_1645;
wire mux_o_1646;
wire mux_o_1647;
wire mux_o_1648;
wire mux_o_1649;
wire mux_o_1650;
wire mux_o_1651;
wire mux_o_1652;
wire mux_o_1653;
wire mux_o_1654;
wire mux_o_1655;
wire mux_o_1656;
wire mux_o_1657;
wire mux_o_1658;
wire mux_o_1659;
wire mux_o_1660;
wire mux_o_1661;
wire mux_o_1662;
wire mux_o_1663;
wire mux_o_1664;
wire mux_o_1665;
wire mux_o_1666;
wire mux_o_1667;
wire mux_o_1668;
wire mux_o_1669;
wire mux_o_1670;
wire mux_o_1671;
wire mux_o_1672;
wire mux_o_1673;
wire mux_o_1674;
wire mux_o_1675;
wire mux_o_1676;
wire mux_o_1677;
wire mux_o_1678;
wire mux_o_1679;
wire mux_o_1680;
wire mux_o_1681;
wire mux_o_1682;
wire mux_o_1683;
wire mux_o_1684;
wire mux_o_1685;
wire mux_o_1686;
wire mux_o_1687;
wire mux_o_1688;
wire mux_o_1689;
wire mux_o_1690;
wire mux_o_1691;
wire mux_o_1692;
wire mux_o_1693;
wire mux_o_1694;
wire mux_o_1695;
wire mux_o_1696;
wire mux_o_1697;
wire mux_o_1698;
wire mux_o_1699;
wire mux_o_1700;
wire mux_o_1701;
wire mux_o_1702;
wire mux_o_1703;
wire mux_o_1704;
wire mux_o_1705;
wire mux_o_1706;
wire mux_o_1707;
wire mux_o_1708;
wire mux_o_1709;
wire mux_o_1710;
wire mux_o_1711;
wire mux_o_1712;
wire mux_o_1713;
wire mux_o_1714;
wire mux_o_1715;
wire mux_o_1716;
wire mux_o_1717;
wire mux_o_1718;
wire mux_o_1719;
wire mux_o_1720;
wire mux_o_1721;
wire mux_o_1722;
wire mux_o_1723;
wire mux_o_1724;
wire mux_o_1725;
wire mux_o_1726;
wire mux_o_1727;
wire mux_o_1728;
wire mux_o_1729;
wire mux_o_1730;
wire mux_o_1731;
wire mux_o_1732;
wire mux_o_1733;
wire mux_o_1734;
wire mux_o_1735;
wire mux_o_1736;
wire mux_o_1737;
wire mux_o_1738;
wire mux_o_1739;
wire mux_o_1740;
wire mux_o_1741;
wire mux_o_1742;
wire mux_o_1743;
wire mux_o_1744;
wire mux_o_1745;
wire mux_o_1746;
wire mux_o_1747;
wire mux_o_1748;
wire mux_o_1749;
wire mux_o_1750;
wire mux_o_1751;
wire mux_o_1752;
wire mux_o_1753;
wire mux_o_1754;
wire mux_o_1755;
wire mux_o_1756;
wire mux_o_1757;
wire mux_o_1758;
wire mux_o_1759;
wire mux_o_1760;
wire mux_o_1761;
wire mux_o_1762;
wire mux_o_1763;
wire mux_o_1764;
wire mux_o_1765;
wire mux_o_1766;
wire mux_o_1767;
wire mux_o_1768;
wire mux_o_1769;
wire mux_o_1770;
wire mux_o_1771;
wire mux_o_1772;
wire mux_o_1773;
wire mux_o_1774;
wire mux_o_1775;
wire mux_o_1776;
wire mux_o_1777;
wire mux_o_1778;
wire mux_o_1779;
wire mux_o_1780;
wire mux_o_1781;
wire mux_o_1782;
wire mux_o_1783;
wire mux_o_1784;
wire mux_o_1785;
wire mux_o_1786;
wire mux_o_1787;
wire mux_o_1788;
wire mux_o_1789;
wire mux_o_1790;
wire mux_o_1791;
wire mux_o_1792;
wire mux_o_1793;
wire mux_o_1794;
wire mux_o_1795;
wire mux_o_1796;
wire mux_o_1797;
wire mux_o_1798;
wire mux_o_1799;
wire mux_o_1800;
wire mux_o_1801;
wire mux_o_1802;
wire mux_o_1803;
wire mux_o_1804;
wire mux_o_1805;
wire mux_o_1806;
wire mux_o_1807;
wire mux_o_1808;
wire mux_o_1809;
wire mux_o_1810;
wire mux_o_1811;
wire mux_o_1812;
wire mux_o_1813;
wire mux_o_1814;
wire mux_o_1815;
wire mux_o_1816;
wire mux_o_1817;
wire mux_o_1818;
wire mux_o_1819;
wire mux_o_1820;
wire mux_o_1821;
wire mux_o_1822;
wire mux_o_1823;
wire mux_o_1824;
wire mux_o_1825;
wire mux_o_1826;
wire mux_o_1827;
wire mux_o_1828;
wire mux_o_1829;
wire mux_o_1830;
wire mux_o_1831;
wire mux_o_1832;
wire mux_o_1833;
wire mux_o_1834;
wire mux_o_1835;
wire mux_o_1836;
wire mux_o_1837;
wire mux_o_1838;
wire mux_o_1839;
wire mux_o_1840;
wire mux_o_1841;
wire mux_o_1842;
wire mux_o_1843;
wire mux_o_1844;
wire mux_o_1845;
wire mux_o_1846;
wire mux_o_1847;
wire mux_o_1848;
wire mux_o_1849;
wire mux_o_1850;
wire mux_o_1851;
wire mux_o_1852;
wire mux_o_1853;
wire mux_o_1854;
wire mux_o_1855;
wire mux_o_1856;
wire mux_o_1857;
wire mux_o_1858;
wire mux_o_1859;
wire mux_o_1860;
wire mux_o_1861;
wire mux_o_1862;
wire mux_o_1863;
wire mux_o_1864;
wire mux_o_1865;
wire mux_o_1866;
wire mux_o_1867;
wire mux_o_1868;
wire mux_o_1869;
wire mux_o_1870;
wire mux_o_1871;
wire mux_o_1872;
wire mux_o_1873;
wire mux_o_1874;
wire mux_o_1875;
wire mux_o_1876;
wire mux_o_1877;
wire mux_o_1878;
wire mux_o_1879;
wire mux_o_1880;
wire mux_o_1881;
wire mux_o_1882;
wire mux_o_1883;
wire mux_o_1884;
wire mux_o_1885;
wire mux_o_1886;
wire mux_o_1887;
wire mux_o_1888;
wire mux_o_1889;
wire mux_o_1890;
wire mux_o_1891;
wire mux_o_1892;
wire mux_o_1893;
wire mux_o_1894;
wire mux_o_1895;
wire mux_o_1896;
wire mux_o_1897;
wire mux_o_1898;
wire mux_o_1899;
wire mux_o_1900;
wire mux_o_1901;
wire mux_o_1902;
wire mux_o_1903;
wire mux_o_1904;
wire mux_o_1905;
wire mux_o_1906;
wire mux_o_1907;
wire mux_o_1908;
wire mux_o_1909;
wire mux_o_1910;
wire mux_o_1911;
wire mux_o_1912;
wire mux_o_1913;
wire mux_o_1914;
wire mux_o_1915;
wire mux_o_1916;
wire mux_o_1917;
wire mux_o_1918;
wire mux_o_1919;
wire mux_o_1920;
wire mux_o_1921;
wire mux_o_1922;
wire mux_o_1923;
wire mux_o_1924;
wire mux_o_1925;
wire mux_o_1926;
wire mux_o_1927;
wire mux_o_1928;
wire mux_o_1929;
wire mux_o_1930;
wire mux_o_1931;
wire mux_o_1932;
wire mux_o_1933;
wire mux_o_1934;
wire mux_o_1935;
wire mux_o_1936;
wire mux_o_1937;
wire mux_o_1938;
wire mux_o_1939;
wire mux_o_1940;
wire mux_o_1941;
wire mux_o_1942;
wire mux_o_1943;
wire mux_o_1944;
wire mux_o_1945;
wire mux_o_1946;
wire mux_o_1947;
wire mux_o_1948;
wire mux_o_1949;
wire mux_o_1950;
wire mux_o_1951;
wire mux_o_1952;
wire mux_o_1953;
wire mux_o_1954;
wire mux_o_1955;
wire mux_o_1956;
wire mux_o_1957;
wire mux_o_1958;
wire mux_o_1959;
wire mux_o_1960;
wire mux_o_1961;
wire mux_o_1962;
wire mux_o_1963;
wire mux_o_1964;
wire mux_o_1965;
wire mux_o_1966;
wire mux_o_1967;
wire mux_o_1968;
wire mux_o_1969;
wire mux_o_1970;
wire mux_o_1971;
wire mux_o_1972;
wire mux_o_1973;
wire mux_o_1974;
wire mux_o_1975;
wire mux_o_1976;
wire mux_o_1977;
wire mux_o_1978;
wire mux_o_1979;
wire mux_o_1980;
wire mux_o_1981;
wire mux_o_1982;
wire mux_o_1983;
wire mux_o_1984;
wire mux_o_1985;
wire mux_o_1986;
wire mux_o_1987;
wire mux_o_1988;
wire mux_o_1989;
wire mux_o_1990;
wire mux_o_1991;
wire mux_o_1992;
wire mux_o_1993;
wire mux_o_1994;
wire mux_o_1995;
wire mux_o_1996;
wire mux_o_1997;
wire mux_o_1998;
wire mux_o_1999;
wire mux_o_2000;
wire mux_o_2001;
wire mux_o_2002;
wire mux_o_2003;
wire mux_o_2004;
wire mux_o_2005;
wire mux_o_2006;
wire mux_o_2007;
wire mux_o_2008;
wire mux_o_2009;
wire mux_o_2010;
wire mux_o_2011;
wire mux_o_2012;
wire mux_o_2013;
wire mux_o_2014;
wire mux_o_2015;
wire mux_o_2016;
wire mux_o_2017;
wire mux_o_2018;
wire mux_o_2019;
wire mux_o_2020;
wire mux_o_2021;
wire mux_o_2022;
wire mux_o_2023;
wire mux_o_2024;
wire mux_o_2025;
wire mux_o_2026;
wire mux_o_2027;
wire mux_o_2028;
wire mux_o_2029;
wire mux_o_2030;
wire mux_o_2031;
wire mux_o_2032;
wire mux_o_2033;
wire mux_o_2034;
wire mux_o_2035;
wire mux_o_2036;
wire mux_o_2037;
wire mux_o_2038;
wire mux_o_2039;
wire mux_o_2040;
wire mux_o_2041;
wire mux_o_2042;
wire mux_o_2043;
wire mux_o_2044;
wire mux_o_2045;
wire mux_o_2046;
wire mux_o_2047;
wire mux_o_2048;
wire mux_o_2049;
wire mux_o_2050;
wire mux_o_2051;
wire mux_o_2052;
wire mux_o_2053;
wire mux_o_2054;
wire mux_o_2055;
wire mux_o_2056;
wire mux_o_2057;
wire mux_o_2058;
wire mux_o_2059;
wire mux_o_2060;
wire mux_o_2061;
wire mux_o_2062;
wire mux_o_2063;
wire mux_o_2064;
wire mux_o_2065;
wire mux_o_2066;
wire mux_o_2067;
wire mux_o_2068;
wire mux_o_2069;
wire mux_o_2070;
wire mux_o_2071;
wire mux_o_2072;
wire mux_o_2073;
wire mux_o_2074;
wire mux_o_2075;
wire mux_o_2076;
wire mux_o_2077;
wire mux_o_2078;
wire mux_o_2079;
wire mux_o_2080;
wire mux_o_2081;
wire mux_o_2082;
wire mux_o_2083;
wire mux_o_2084;
wire mux_o_2085;
wire mux_o_2086;
wire mux_o_2087;
wire mux_o_2088;
wire mux_o_2089;
wire mux_o_2090;
wire mux_o_2091;
wire mux_o_2092;
wire mux_o_2093;
wire mux_o_2094;
wire mux_o_2095;
wire mux_o_2096;
wire mux_o_2097;
wire mux_o_2098;
wire mux_o_2099;
wire mux_o_2100;
wire mux_o_2101;
wire mux_o_2102;
wire mux_o_2103;
wire mux_o_2104;
wire mux_o_2105;
wire mux_o_2106;
wire mux_o_2107;
wire mux_o_2108;
wire mux_o_2109;
wire mux_o_2110;
wire mux_o_2111;
wire mux_o_2112;
wire mux_o_2113;
wire mux_o_2114;
wire mux_o_2115;
wire mux_o_2116;
wire mux_o_2117;
wire mux_o_2118;
wire mux_o_2119;
wire mux_o_2120;
wire mux_o_2121;
wire mux_o_2122;
wire mux_o_2123;
wire mux_o_2124;
wire mux_o_2125;
wire mux_o_2126;
wire mux_o_2127;
wire mux_o_2128;
wire mux_o_2129;
wire mux_o_2130;
wire mux_o_2131;
wire mux_o_2132;
wire mux_o_2133;
wire mux_o_2134;
wire mux_o_2135;
wire mux_o_2136;
wire mux_o_2137;
wire mux_o_2138;
wire mux_o_2139;
wire mux_o_2140;
wire mux_o_2141;
wire mux_o_2142;
wire mux_o_2143;
wire mux_o_2144;
wire mux_o_2145;
wire mux_o_2146;
wire mux_o_2147;
wire mux_o_2148;
wire mux_o_2149;
wire mux_o_2150;
wire mux_o_2151;
wire mux_o_2152;
wire mux_o_2153;
wire mux_o_2154;
wire mux_o_2155;
wire mux_o_2156;
wire mux_o_2157;
wire mux_o_2158;
wire mux_o_2159;
wire mux_o_2160;
wire mux_o_2161;
wire mux_o_2162;
wire mux_o_2163;
wire mux_o_2164;
wire mux_o_2165;
wire mux_o_2166;
wire mux_o_2167;
wire mux_o_2168;
wire mux_o_2169;
wire mux_o_2170;
wire mux_o_2171;
wire mux_o_2172;
wire mux_o_2173;
wire mux_o_2174;
wire mux_o_2175;
wire mux_o_2176;
wire mux_o_2177;
wire mux_o_2178;
wire mux_o_2179;
wire mux_o_2180;
wire mux_o_2181;
wire mux_o_2182;
wire mux_o_2183;
wire mux_o_2184;
wire mux_o_2185;
wire mux_o_2186;
wire mux_o_2187;
wire mux_o_2188;
wire mux_o_2189;
wire mux_o_2190;
wire mux_o_2191;
wire mux_o_2192;
wire mux_o_2193;
wire mux_o_2194;
wire mux_o_2195;
wire mux_o_2196;
wire mux_o_2197;
wire mux_o_2198;
wire mux_o_2199;
wire mux_o_2200;
wire mux_o_2201;
wire mux_o_2202;
wire mux_o_2203;
wire mux_o_2204;
wire mux_o_2205;
wire mux_o_2206;
wire mux_o_2207;
wire mux_o_2208;
wire mux_o_2209;
wire mux_o_2210;
wire mux_o_2211;
wire mux_o_2212;
wire mux_o_2213;
wire mux_o_2214;
wire mux_o_2215;
wire mux_o_2216;
wire mux_o_2217;
wire mux_o_2218;
wire mux_o_2219;
wire mux_o_2220;
wire mux_o_2221;
wire mux_o_2222;
wire mux_o_2223;
wire mux_o_2224;
wire mux_o_2225;
wire mux_o_2226;
wire mux_o_2227;
wire mux_o_2228;
wire mux_o_2229;
wire mux_o_2230;
wire mux_o_2231;
wire mux_o_2232;
wire mux_o_2233;
wire mux_o_2234;
wire mux_o_2235;
wire mux_o_2236;
wire mux_o_2237;
wire mux_o_2238;
wire mux_o_2239;
wire mux_o_2240;
wire mux_o_2241;
wire mux_o_2242;
wire mux_o_2243;
wire mux_o_2244;
wire mux_o_2245;
wire mux_o_2246;
wire mux_o_2247;
wire mux_o_2248;
wire mux_o_2249;
wire mux_o_2250;
wire mux_o_2251;
wire mux_o_2252;
wire mux_o_2253;
wire mux_o_2254;
wire mux_o_2255;
wire mux_o_2256;
wire mux_o_2257;
wire mux_o_2258;
wire mux_o_2259;
wire mux_o_2260;
wire mux_o_2261;
wire mux_o_2262;
wire mux_o_2263;
wire mux_o_2264;
wire mux_o_2265;
wire mux_o_2266;
wire mux_o_2267;
wire mux_o_2268;
wire mux_o_2269;
wire mux_o_2270;
wire mux_o_2271;
wire mux_o_2272;
wire mux_o_2273;
wire mux_o_2274;
wire mux_o_2275;
wire mux_o_2276;
wire mux_o_2277;
wire mux_o_2278;
wire mux_o_2279;
wire mux_o_2280;
wire mux_o_2281;
wire mux_o_2282;
wire mux_o_2283;
wire mux_o_2284;
wire mux_o_2285;
wire mux_o_2286;
wire mux_o_2287;
wire mux_o_2288;
wire mux_o_2289;
wire mux_o_2290;
wire mux_o_2291;
wire mux_o_2292;
wire mux_o_2293;
wire mux_o_2294;
wire mux_o_2295;
wire mux_o_2296;
wire mux_o_2297;
wire mux_o_2298;
wire mux_o_2299;
wire mux_o_2300;
wire mux_o_2301;
wire mux_o_2302;
wire mux_o_2303;
wire mux_o_2304;
wire mux_o_2305;
wire mux_o_2306;
wire mux_o_2307;
wire mux_o_2308;
wire mux_o_2309;
wire mux_o_2310;
wire mux_o_2311;
wire mux_o_2312;
wire mux_o_2313;
wire mux_o_2314;
wire mux_o_2315;
wire mux_o_2316;
wire mux_o_2317;
wire mux_o_2318;
wire mux_o_2319;
wire mux_o_2320;
wire mux_o_2321;
wire mux_o_2322;
wire mux_o_2323;
wire mux_o_2324;
wire mux_o_2325;
wire mux_o_2326;
wire mux_o_2327;
wire mux_o_2328;
wire mux_o_2329;
wire mux_o_2330;
wire mux_o_2331;
wire mux_o_2332;
wire mux_o_2333;
wire mux_o_2334;
wire mux_o_2335;
wire mux_o_2336;
wire mux_o_2337;
wire mux_o_2338;
wire mux_o_2339;
wire mux_o_2340;
wire mux_o_2341;
wire mux_o_2342;
wire mux_o_2343;
wire mux_o_2344;
wire mux_o_2345;
wire mux_o_2346;
wire mux_o_2347;
wire mux_o_2348;
wire mux_o_2349;
wire mux_o_2350;
wire mux_o_2351;
wire mux_o_2352;
wire mux_o_2353;
wire mux_o_2354;
wire mux_o_2355;
wire mux_o_2356;
wire mux_o_2357;
wire mux_o_2358;
wire mux_o_2359;
wire mux_o_2360;
wire mux_o_2361;
wire mux_o_2362;
wire mux_o_2363;
wire mux_o_2364;
wire mux_o_2365;
wire mux_o_2366;
wire mux_o_2367;
wire mux_o_2368;
wire mux_o_2369;
wire mux_o_2370;
wire mux_o_2371;
wire mux_o_2372;
wire mux_o_2373;
wire mux_o_2374;
wire mux_o_2375;
wire mux_o_2376;
wire mux_o_2377;
wire mux_o_2378;
wire mux_o_2379;
wire mux_o_2380;
wire mux_o_2381;
wire mux_o_2382;
wire mux_o_2383;
wire mux_o_2384;
wire mux_o_2385;
wire mux_o_2386;
wire mux_o_2387;
wire mux_o_2388;
wire mux_o_2389;
wire mux_o_2390;
wire mux_o_2392;
wire mux_o_2393;
wire mux_o_2394;
wire mux_o_2395;
wire mux_o_2396;
wire mux_o_2397;
wire mux_o_2399;
wire mux_o_2400;
wire mux_o_2401;
wire mux_o_2403;
wire mux_o_2404;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

INV inv_inst_0 (.I(ad[4]), .O(ad4_inv));

INV inv_inst_1 (.I(ad[5]), .O(ad5_inv));

INV inv_inst_2 (.I(ad[6]), .O(ad6_inv));

INV inv_inst_3 (.I(ad[7]), .O(ad7_inv));

INV inv_inst_4 (.I(ad[8]), .O(ad8_inv));

INV inv_inst_5 (.I(ad[9]), .O(ad9_inv));

INV inv_inst_6 (.I(ad[10]), .O(ad10_inv));

INV inv_inst_7 (.I(ad[11]), .O(ad11_inv));

INV inv_inst_8 (.I(ad[12]), .O(ad12_inv));

INV inv_inst_9 (.I(ad[13]), .O(ad13_inv));

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_0.INIT = 16'h8000;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1.INIT = 16'h8000;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_2.INIT = 16'h8000;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(lut_f_0),
  .I1(lut_f_1),
  .I2(lut_f_2),
  .I3(gw_vcc)
);
defparam lut_inst_3.INIT = 16'h8000;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_4.INIT = 16'h8000;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_5.INIT = 16'h8000;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_6.INIT = 16'h8000;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(lut_f_4),
  .I1(lut_f_5),
  .I2(lut_f_6),
  .I3(gw_vcc)
);
defparam lut_inst_7.INIT = 16'h8000;
LUT4 lut_inst_8 (
  .F(lut_f_8),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_8.INIT = 16'h8000;
LUT4 lut_inst_9 (
  .F(lut_f_9),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_9.INIT = 16'h8000;
LUT4 lut_inst_10 (
  .F(lut_f_10),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_10.INIT = 16'h8000;
LUT4 lut_inst_11 (
  .F(lut_f_11),
  .I0(lut_f_8),
  .I1(lut_f_9),
  .I2(lut_f_10),
  .I3(gw_vcc)
);
defparam lut_inst_11.INIT = 16'h8000;
LUT4 lut_inst_12 (
  .F(lut_f_12),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_12.INIT = 16'h8000;
LUT4 lut_inst_13 (
  .F(lut_f_13),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_13.INIT = 16'h8000;
LUT4 lut_inst_14 (
  .F(lut_f_14),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_14.INIT = 16'h8000;
LUT4 lut_inst_15 (
  .F(lut_f_15),
  .I0(lut_f_12),
  .I1(lut_f_13),
  .I2(lut_f_14),
  .I3(gw_vcc)
);
defparam lut_inst_15.INIT = 16'h8000;
LUT4 lut_inst_16 (
  .F(lut_f_16),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_16.INIT = 16'h8000;
LUT4 lut_inst_17 (
  .F(lut_f_17),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_17.INIT = 16'h8000;
LUT4 lut_inst_18 (
  .F(lut_f_18),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_18.INIT = 16'h8000;
LUT4 lut_inst_19 (
  .F(lut_f_19),
  .I0(lut_f_16),
  .I1(lut_f_17),
  .I2(lut_f_18),
  .I3(gw_vcc)
);
defparam lut_inst_19.INIT = 16'h8000;
LUT4 lut_inst_20 (
  .F(lut_f_20),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_20.INIT = 16'h8000;
LUT4 lut_inst_21 (
  .F(lut_f_21),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_21.INIT = 16'h8000;
LUT4 lut_inst_22 (
  .F(lut_f_22),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_22.INIT = 16'h8000;
LUT4 lut_inst_23 (
  .F(lut_f_23),
  .I0(lut_f_20),
  .I1(lut_f_21),
  .I2(lut_f_22),
  .I3(gw_vcc)
);
defparam lut_inst_23.INIT = 16'h8000;
LUT4 lut_inst_24 (
  .F(lut_f_24),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_24.INIT = 16'h8000;
LUT4 lut_inst_25 (
  .F(lut_f_25),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_25.INIT = 16'h8000;
LUT4 lut_inst_26 (
  .F(lut_f_26),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_26.INIT = 16'h8000;
LUT4 lut_inst_27 (
  .F(lut_f_27),
  .I0(lut_f_24),
  .I1(lut_f_25),
  .I2(lut_f_26),
  .I3(gw_vcc)
);
defparam lut_inst_27.INIT = 16'h8000;
LUT4 lut_inst_28 (
  .F(lut_f_28),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_28.INIT = 16'h8000;
LUT4 lut_inst_29 (
  .F(lut_f_29),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_29.INIT = 16'h8000;
LUT4 lut_inst_30 (
  .F(lut_f_30),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_30.INIT = 16'h8000;
LUT4 lut_inst_31 (
  .F(lut_f_31),
  .I0(lut_f_28),
  .I1(lut_f_29),
  .I2(lut_f_30),
  .I3(gw_vcc)
);
defparam lut_inst_31.INIT = 16'h8000;
LUT4 lut_inst_32 (
  .F(lut_f_32),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_32.INIT = 16'h8000;
LUT4 lut_inst_33 (
  .F(lut_f_33),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_33.INIT = 16'h8000;
LUT4 lut_inst_34 (
  .F(lut_f_34),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_34.INIT = 16'h8000;
LUT4 lut_inst_35 (
  .F(lut_f_35),
  .I0(lut_f_32),
  .I1(lut_f_33),
  .I2(lut_f_34),
  .I3(gw_vcc)
);
defparam lut_inst_35.INIT = 16'h8000;
LUT4 lut_inst_36 (
  .F(lut_f_36),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_36.INIT = 16'h8000;
LUT4 lut_inst_37 (
  .F(lut_f_37),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_37.INIT = 16'h8000;
LUT4 lut_inst_38 (
  .F(lut_f_38),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_38.INIT = 16'h8000;
LUT4 lut_inst_39 (
  .F(lut_f_39),
  .I0(lut_f_36),
  .I1(lut_f_37),
  .I2(lut_f_38),
  .I3(gw_vcc)
);
defparam lut_inst_39.INIT = 16'h8000;
LUT4 lut_inst_40 (
  .F(lut_f_40),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_40.INIT = 16'h8000;
LUT4 lut_inst_41 (
  .F(lut_f_41),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_41.INIT = 16'h8000;
LUT4 lut_inst_42 (
  .F(lut_f_42),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_42.INIT = 16'h8000;
LUT4 lut_inst_43 (
  .F(lut_f_43),
  .I0(lut_f_40),
  .I1(lut_f_41),
  .I2(lut_f_42),
  .I3(gw_vcc)
);
defparam lut_inst_43.INIT = 16'h8000;
LUT4 lut_inst_44 (
  .F(lut_f_44),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_44.INIT = 16'h8000;
LUT4 lut_inst_45 (
  .F(lut_f_45),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_45.INIT = 16'h8000;
LUT4 lut_inst_46 (
  .F(lut_f_46),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_46.INIT = 16'h8000;
LUT4 lut_inst_47 (
  .F(lut_f_47),
  .I0(lut_f_44),
  .I1(lut_f_45),
  .I2(lut_f_46),
  .I3(gw_vcc)
);
defparam lut_inst_47.INIT = 16'h8000;
LUT4 lut_inst_48 (
  .F(lut_f_48),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_48.INIT = 16'h8000;
LUT4 lut_inst_49 (
  .F(lut_f_49),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_49.INIT = 16'h8000;
LUT4 lut_inst_50 (
  .F(lut_f_50),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_50.INIT = 16'h8000;
LUT4 lut_inst_51 (
  .F(lut_f_51),
  .I0(lut_f_48),
  .I1(lut_f_49),
  .I2(lut_f_50),
  .I3(gw_vcc)
);
defparam lut_inst_51.INIT = 16'h8000;
LUT4 lut_inst_52 (
  .F(lut_f_52),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_52.INIT = 16'h8000;
LUT4 lut_inst_53 (
  .F(lut_f_53),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_53.INIT = 16'h8000;
LUT4 lut_inst_54 (
  .F(lut_f_54),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_54.INIT = 16'h8000;
LUT4 lut_inst_55 (
  .F(lut_f_55),
  .I0(lut_f_52),
  .I1(lut_f_53),
  .I2(lut_f_54),
  .I3(gw_vcc)
);
defparam lut_inst_55.INIT = 16'h8000;
LUT4 lut_inst_56 (
  .F(lut_f_56),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_56.INIT = 16'h8000;
LUT4 lut_inst_57 (
  .F(lut_f_57),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_57.INIT = 16'h8000;
LUT4 lut_inst_58 (
  .F(lut_f_58),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_58.INIT = 16'h8000;
LUT4 lut_inst_59 (
  .F(lut_f_59),
  .I0(lut_f_56),
  .I1(lut_f_57),
  .I2(lut_f_58),
  .I3(gw_vcc)
);
defparam lut_inst_59.INIT = 16'h8000;
LUT4 lut_inst_60 (
  .F(lut_f_60),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_60.INIT = 16'h8000;
LUT4 lut_inst_61 (
  .F(lut_f_61),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_61.INIT = 16'h8000;
LUT4 lut_inst_62 (
  .F(lut_f_62),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_62.INIT = 16'h8000;
LUT4 lut_inst_63 (
  .F(lut_f_63),
  .I0(lut_f_60),
  .I1(lut_f_61),
  .I2(lut_f_62),
  .I3(gw_vcc)
);
defparam lut_inst_63.INIT = 16'h8000;
LUT4 lut_inst_64 (
  .F(lut_f_64),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_64.INIT = 16'h8000;
LUT4 lut_inst_65 (
  .F(lut_f_65),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_65.INIT = 16'h8000;
LUT4 lut_inst_66 (
  .F(lut_f_66),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_66.INIT = 16'h8000;
LUT4 lut_inst_67 (
  .F(lut_f_67),
  .I0(lut_f_64),
  .I1(lut_f_65),
  .I2(lut_f_66),
  .I3(gw_vcc)
);
defparam lut_inst_67.INIT = 16'h8000;
LUT4 lut_inst_68 (
  .F(lut_f_68),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_68.INIT = 16'h8000;
LUT4 lut_inst_69 (
  .F(lut_f_69),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_69.INIT = 16'h8000;
LUT4 lut_inst_70 (
  .F(lut_f_70),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_70.INIT = 16'h8000;
LUT4 lut_inst_71 (
  .F(lut_f_71),
  .I0(lut_f_68),
  .I1(lut_f_69),
  .I2(lut_f_70),
  .I3(gw_vcc)
);
defparam lut_inst_71.INIT = 16'h8000;
LUT4 lut_inst_72 (
  .F(lut_f_72),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_72.INIT = 16'h8000;
LUT4 lut_inst_73 (
  .F(lut_f_73),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_73.INIT = 16'h8000;
LUT4 lut_inst_74 (
  .F(lut_f_74),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_74.INIT = 16'h8000;
LUT4 lut_inst_75 (
  .F(lut_f_75),
  .I0(lut_f_72),
  .I1(lut_f_73),
  .I2(lut_f_74),
  .I3(gw_vcc)
);
defparam lut_inst_75.INIT = 16'h8000;
LUT4 lut_inst_76 (
  .F(lut_f_76),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_76.INIT = 16'h8000;
LUT4 lut_inst_77 (
  .F(lut_f_77),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_77.INIT = 16'h8000;
LUT4 lut_inst_78 (
  .F(lut_f_78),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_78.INIT = 16'h8000;
LUT4 lut_inst_79 (
  .F(lut_f_79),
  .I0(lut_f_76),
  .I1(lut_f_77),
  .I2(lut_f_78),
  .I3(gw_vcc)
);
defparam lut_inst_79.INIT = 16'h8000;
LUT4 lut_inst_80 (
  .F(lut_f_80),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_80.INIT = 16'h8000;
LUT4 lut_inst_81 (
  .F(lut_f_81),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_81.INIT = 16'h8000;
LUT4 lut_inst_82 (
  .F(lut_f_82),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_82.INIT = 16'h8000;
LUT4 lut_inst_83 (
  .F(lut_f_83),
  .I0(lut_f_80),
  .I1(lut_f_81),
  .I2(lut_f_82),
  .I3(gw_vcc)
);
defparam lut_inst_83.INIT = 16'h8000;
LUT4 lut_inst_84 (
  .F(lut_f_84),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_84.INIT = 16'h8000;
LUT4 lut_inst_85 (
  .F(lut_f_85),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_85.INIT = 16'h8000;
LUT4 lut_inst_86 (
  .F(lut_f_86),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_86.INIT = 16'h8000;
LUT4 lut_inst_87 (
  .F(lut_f_87),
  .I0(lut_f_84),
  .I1(lut_f_85),
  .I2(lut_f_86),
  .I3(gw_vcc)
);
defparam lut_inst_87.INIT = 16'h8000;
LUT4 lut_inst_88 (
  .F(lut_f_88),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_88.INIT = 16'h8000;
LUT4 lut_inst_89 (
  .F(lut_f_89),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_89.INIT = 16'h8000;
LUT4 lut_inst_90 (
  .F(lut_f_90),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_90.INIT = 16'h8000;
LUT4 lut_inst_91 (
  .F(lut_f_91),
  .I0(lut_f_88),
  .I1(lut_f_89),
  .I2(lut_f_90),
  .I3(gw_vcc)
);
defparam lut_inst_91.INIT = 16'h8000;
LUT4 lut_inst_92 (
  .F(lut_f_92),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_92.INIT = 16'h8000;
LUT4 lut_inst_93 (
  .F(lut_f_93),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_93.INIT = 16'h8000;
LUT4 lut_inst_94 (
  .F(lut_f_94),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_94.INIT = 16'h8000;
LUT4 lut_inst_95 (
  .F(lut_f_95),
  .I0(lut_f_92),
  .I1(lut_f_93),
  .I2(lut_f_94),
  .I3(gw_vcc)
);
defparam lut_inst_95.INIT = 16'h8000;
LUT4 lut_inst_96 (
  .F(lut_f_96),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_96.INIT = 16'h8000;
LUT4 lut_inst_97 (
  .F(lut_f_97),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_97.INIT = 16'h8000;
LUT4 lut_inst_98 (
  .F(lut_f_98),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_98.INIT = 16'h8000;
LUT4 lut_inst_99 (
  .F(lut_f_99),
  .I0(lut_f_96),
  .I1(lut_f_97),
  .I2(lut_f_98),
  .I3(gw_vcc)
);
defparam lut_inst_99.INIT = 16'h8000;
LUT4 lut_inst_100 (
  .F(lut_f_100),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_100.INIT = 16'h8000;
LUT4 lut_inst_101 (
  .F(lut_f_101),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_101.INIT = 16'h8000;
LUT4 lut_inst_102 (
  .F(lut_f_102),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_102.INIT = 16'h8000;
LUT4 lut_inst_103 (
  .F(lut_f_103),
  .I0(lut_f_100),
  .I1(lut_f_101),
  .I2(lut_f_102),
  .I3(gw_vcc)
);
defparam lut_inst_103.INIT = 16'h8000;
LUT4 lut_inst_104 (
  .F(lut_f_104),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_104.INIT = 16'h8000;
LUT4 lut_inst_105 (
  .F(lut_f_105),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_105.INIT = 16'h8000;
LUT4 lut_inst_106 (
  .F(lut_f_106),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_106.INIT = 16'h8000;
LUT4 lut_inst_107 (
  .F(lut_f_107),
  .I0(lut_f_104),
  .I1(lut_f_105),
  .I2(lut_f_106),
  .I3(gw_vcc)
);
defparam lut_inst_107.INIT = 16'h8000;
LUT4 lut_inst_108 (
  .F(lut_f_108),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_108.INIT = 16'h8000;
LUT4 lut_inst_109 (
  .F(lut_f_109),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_109.INIT = 16'h8000;
LUT4 lut_inst_110 (
  .F(lut_f_110),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_110.INIT = 16'h8000;
LUT4 lut_inst_111 (
  .F(lut_f_111),
  .I0(lut_f_108),
  .I1(lut_f_109),
  .I2(lut_f_110),
  .I3(gw_vcc)
);
defparam lut_inst_111.INIT = 16'h8000;
LUT4 lut_inst_112 (
  .F(lut_f_112),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_112.INIT = 16'h8000;
LUT4 lut_inst_113 (
  .F(lut_f_113),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_113.INIT = 16'h8000;
LUT4 lut_inst_114 (
  .F(lut_f_114),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_114.INIT = 16'h8000;
LUT4 lut_inst_115 (
  .F(lut_f_115),
  .I0(lut_f_112),
  .I1(lut_f_113),
  .I2(lut_f_114),
  .I3(gw_vcc)
);
defparam lut_inst_115.INIT = 16'h8000;
LUT4 lut_inst_116 (
  .F(lut_f_116),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_116.INIT = 16'h8000;
LUT4 lut_inst_117 (
  .F(lut_f_117),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_117.INIT = 16'h8000;
LUT4 lut_inst_118 (
  .F(lut_f_118),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_118.INIT = 16'h8000;
LUT4 lut_inst_119 (
  .F(lut_f_119),
  .I0(lut_f_116),
  .I1(lut_f_117),
  .I2(lut_f_118),
  .I3(gw_vcc)
);
defparam lut_inst_119.INIT = 16'h8000;
LUT4 lut_inst_120 (
  .F(lut_f_120),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_120.INIT = 16'h8000;
LUT4 lut_inst_121 (
  .F(lut_f_121),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_121.INIT = 16'h8000;
LUT4 lut_inst_122 (
  .F(lut_f_122),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_122.INIT = 16'h8000;
LUT4 lut_inst_123 (
  .F(lut_f_123),
  .I0(lut_f_120),
  .I1(lut_f_121),
  .I2(lut_f_122),
  .I3(gw_vcc)
);
defparam lut_inst_123.INIT = 16'h8000;
LUT4 lut_inst_124 (
  .F(lut_f_124),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_124.INIT = 16'h8000;
LUT4 lut_inst_125 (
  .F(lut_f_125),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_125.INIT = 16'h8000;
LUT4 lut_inst_126 (
  .F(lut_f_126),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_126.INIT = 16'h8000;
LUT4 lut_inst_127 (
  .F(lut_f_127),
  .I0(lut_f_124),
  .I1(lut_f_125),
  .I2(lut_f_126),
  .I3(gw_vcc)
);
defparam lut_inst_127.INIT = 16'h8000;
LUT4 lut_inst_128 (
  .F(lut_f_128),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_128.INIT = 16'h8000;
LUT4 lut_inst_129 (
  .F(lut_f_129),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_129.INIT = 16'h8000;
LUT4 lut_inst_130 (
  .F(lut_f_130),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_130.INIT = 16'h8000;
LUT4 lut_inst_131 (
  .F(lut_f_131),
  .I0(lut_f_128),
  .I1(lut_f_129),
  .I2(lut_f_130),
  .I3(gw_vcc)
);
defparam lut_inst_131.INIT = 16'h8000;
LUT4 lut_inst_132 (
  .F(lut_f_132),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_132.INIT = 16'h8000;
LUT4 lut_inst_133 (
  .F(lut_f_133),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_133.INIT = 16'h8000;
LUT4 lut_inst_134 (
  .F(lut_f_134),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_134.INIT = 16'h8000;
LUT4 lut_inst_135 (
  .F(lut_f_135),
  .I0(lut_f_132),
  .I1(lut_f_133),
  .I2(lut_f_134),
  .I3(gw_vcc)
);
defparam lut_inst_135.INIT = 16'h8000;
LUT4 lut_inst_136 (
  .F(lut_f_136),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_136.INIT = 16'h8000;
LUT4 lut_inst_137 (
  .F(lut_f_137),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_137.INIT = 16'h8000;
LUT4 lut_inst_138 (
  .F(lut_f_138),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_138.INIT = 16'h8000;
LUT4 lut_inst_139 (
  .F(lut_f_139),
  .I0(lut_f_136),
  .I1(lut_f_137),
  .I2(lut_f_138),
  .I3(gw_vcc)
);
defparam lut_inst_139.INIT = 16'h8000;
LUT4 lut_inst_140 (
  .F(lut_f_140),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_140.INIT = 16'h8000;
LUT4 lut_inst_141 (
  .F(lut_f_141),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_141.INIT = 16'h8000;
LUT4 lut_inst_142 (
  .F(lut_f_142),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_142.INIT = 16'h8000;
LUT4 lut_inst_143 (
  .F(lut_f_143),
  .I0(lut_f_140),
  .I1(lut_f_141),
  .I2(lut_f_142),
  .I3(gw_vcc)
);
defparam lut_inst_143.INIT = 16'h8000;
LUT4 lut_inst_144 (
  .F(lut_f_144),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_144.INIT = 16'h8000;
LUT4 lut_inst_145 (
  .F(lut_f_145),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_145.INIT = 16'h8000;
LUT4 lut_inst_146 (
  .F(lut_f_146),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_146.INIT = 16'h8000;
LUT4 lut_inst_147 (
  .F(lut_f_147),
  .I0(lut_f_144),
  .I1(lut_f_145),
  .I2(lut_f_146),
  .I3(gw_vcc)
);
defparam lut_inst_147.INIT = 16'h8000;
LUT4 lut_inst_148 (
  .F(lut_f_148),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_148.INIT = 16'h8000;
LUT4 lut_inst_149 (
  .F(lut_f_149),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_149.INIT = 16'h8000;
LUT4 lut_inst_150 (
  .F(lut_f_150),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_150.INIT = 16'h8000;
LUT4 lut_inst_151 (
  .F(lut_f_151),
  .I0(lut_f_148),
  .I1(lut_f_149),
  .I2(lut_f_150),
  .I3(gw_vcc)
);
defparam lut_inst_151.INIT = 16'h8000;
LUT4 lut_inst_152 (
  .F(lut_f_152),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_152.INIT = 16'h8000;
LUT4 lut_inst_153 (
  .F(lut_f_153),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_153.INIT = 16'h8000;
LUT4 lut_inst_154 (
  .F(lut_f_154),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_154.INIT = 16'h8000;
LUT4 lut_inst_155 (
  .F(lut_f_155),
  .I0(lut_f_152),
  .I1(lut_f_153),
  .I2(lut_f_154),
  .I3(gw_vcc)
);
defparam lut_inst_155.INIT = 16'h8000;
LUT4 lut_inst_156 (
  .F(lut_f_156),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_156.INIT = 16'h8000;
LUT4 lut_inst_157 (
  .F(lut_f_157),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_157.INIT = 16'h8000;
LUT4 lut_inst_158 (
  .F(lut_f_158),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_158.INIT = 16'h8000;
LUT4 lut_inst_159 (
  .F(lut_f_159),
  .I0(lut_f_156),
  .I1(lut_f_157),
  .I2(lut_f_158),
  .I3(gw_vcc)
);
defparam lut_inst_159.INIT = 16'h8000;
LUT4 lut_inst_160 (
  .F(lut_f_160),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_160.INIT = 16'h8000;
LUT4 lut_inst_161 (
  .F(lut_f_161),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_161.INIT = 16'h8000;
LUT4 lut_inst_162 (
  .F(lut_f_162),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_162.INIT = 16'h8000;
LUT4 lut_inst_163 (
  .F(lut_f_163),
  .I0(lut_f_160),
  .I1(lut_f_161),
  .I2(lut_f_162),
  .I3(gw_vcc)
);
defparam lut_inst_163.INIT = 16'h8000;
LUT4 lut_inst_164 (
  .F(lut_f_164),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_164.INIT = 16'h8000;
LUT4 lut_inst_165 (
  .F(lut_f_165),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_165.INIT = 16'h8000;
LUT4 lut_inst_166 (
  .F(lut_f_166),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_166.INIT = 16'h8000;
LUT4 lut_inst_167 (
  .F(lut_f_167),
  .I0(lut_f_164),
  .I1(lut_f_165),
  .I2(lut_f_166),
  .I3(gw_vcc)
);
defparam lut_inst_167.INIT = 16'h8000;
LUT4 lut_inst_168 (
  .F(lut_f_168),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_168.INIT = 16'h8000;
LUT4 lut_inst_169 (
  .F(lut_f_169),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_169.INIT = 16'h8000;
LUT4 lut_inst_170 (
  .F(lut_f_170),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_170.INIT = 16'h8000;
LUT4 lut_inst_171 (
  .F(lut_f_171),
  .I0(lut_f_168),
  .I1(lut_f_169),
  .I2(lut_f_170),
  .I3(gw_vcc)
);
defparam lut_inst_171.INIT = 16'h8000;
LUT4 lut_inst_172 (
  .F(lut_f_172),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_172.INIT = 16'h8000;
LUT4 lut_inst_173 (
  .F(lut_f_173),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_173.INIT = 16'h8000;
LUT4 lut_inst_174 (
  .F(lut_f_174),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_174.INIT = 16'h8000;
LUT4 lut_inst_175 (
  .F(lut_f_175),
  .I0(lut_f_172),
  .I1(lut_f_173),
  .I2(lut_f_174),
  .I3(gw_vcc)
);
defparam lut_inst_175.INIT = 16'h8000;
LUT4 lut_inst_176 (
  .F(lut_f_176),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_176.INIT = 16'h8000;
LUT4 lut_inst_177 (
  .F(lut_f_177),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_177.INIT = 16'h8000;
LUT4 lut_inst_178 (
  .F(lut_f_178),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_178.INIT = 16'h8000;
LUT4 lut_inst_179 (
  .F(lut_f_179),
  .I0(lut_f_176),
  .I1(lut_f_177),
  .I2(lut_f_178),
  .I3(gw_vcc)
);
defparam lut_inst_179.INIT = 16'h8000;
LUT4 lut_inst_180 (
  .F(lut_f_180),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_180.INIT = 16'h8000;
LUT4 lut_inst_181 (
  .F(lut_f_181),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_181.INIT = 16'h8000;
LUT4 lut_inst_182 (
  .F(lut_f_182),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_182.INIT = 16'h8000;
LUT4 lut_inst_183 (
  .F(lut_f_183),
  .I0(lut_f_180),
  .I1(lut_f_181),
  .I2(lut_f_182),
  .I3(gw_vcc)
);
defparam lut_inst_183.INIT = 16'h8000;
LUT4 lut_inst_184 (
  .F(lut_f_184),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_184.INIT = 16'h8000;
LUT4 lut_inst_185 (
  .F(lut_f_185),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_185.INIT = 16'h8000;
LUT4 lut_inst_186 (
  .F(lut_f_186),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_186.INIT = 16'h8000;
LUT4 lut_inst_187 (
  .F(lut_f_187),
  .I0(lut_f_184),
  .I1(lut_f_185),
  .I2(lut_f_186),
  .I3(gw_vcc)
);
defparam lut_inst_187.INIT = 16'h8000;
LUT4 lut_inst_188 (
  .F(lut_f_188),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_188.INIT = 16'h8000;
LUT4 lut_inst_189 (
  .F(lut_f_189),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_189.INIT = 16'h8000;
LUT4 lut_inst_190 (
  .F(lut_f_190),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_190.INIT = 16'h8000;
LUT4 lut_inst_191 (
  .F(lut_f_191),
  .I0(lut_f_188),
  .I1(lut_f_189),
  .I2(lut_f_190),
  .I3(gw_vcc)
);
defparam lut_inst_191.INIT = 16'h8000;
LUT4 lut_inst_192 (
  .F(lut_f_192),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_192.INIT = 16'h8000;
LUT4 lut_inst_193 (
  .F(lut_f_193),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_193.INIT = 16'h8000;
LUT4 lut_inst_194 (
  .F(lut_f_194),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_194.INIT = 16'h8000;
LUT4 lut_inst_195 (
  .F(lut_f_195),
  .I0(lut_f_192),
  .I1(lut_f_193),
  .I2(lut_f_194),
  .I3(gw_vcc)
);
defparam lut_inst_195.INIT = 16'h8000;
LUT4 lut_inst_196 (
  .F(lut_f_196),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_196.INIT = 16'h8000;
LUT4 lut_inst_197 (
  .F(lut_f_197),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_197.INIT = 16'h8000;
LUT4 lut_inst_198 (
  .F(lut_f_198),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_198.INIT = 16'h8000;
LUT4 lut_inst_199 (
  .F(lut_f_199),
  .I0(lut_f_196),
  .I1(lut_f_197),
  .I2(lut_f_198),
  .I3(gw_vcc)
);
defparam lut_inst_199.INIT = 16'h8000;
LUT4 lut_inst_200 (
  .F(lut_f_200),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_200.INIT = 16'h8000;
LUT4 lut_inst_201 (
  .F(lut_f_201),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_201.INIT = 16'h8000;
LUT4 lut_inst_202 (
  .F(lut_f_202),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_202.INIT = 16'h8000;
LUT4 lut_inst_203 (
  .F(lut_f_203),
  .I0(lut_f_200),
  .I1(lut_f_201),
  .I2(lut_f_202),
  .I3(gw_vcc)
);
defparam lut_inst_203.INIT = 16'h8000;
LUT4 lut_inst_204 (
  .F(lut_f_204),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_204.INIT = 16'h8000;
LUT4 lut_inst_205 (
  .F(lut_f_205),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_205.INIT = 16'h8000;
LUT4 lut_inst_206 (
  .F(lut_f_206),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_206.INIT = 16'h8000;
LUT4 lut_inst_207 (
  .F(lut_f_207),
  .I0(lut_f_204),
  .I1(lut_f_205),
  .I2(lut_f_206),
  .I3(gw_vcc)
);
defparam lut_inst_207.INIT = 16'h8000;
LUT4 lut_inst_208 (
  .F(lut_f_208),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_208.INIT = 16'h8000;
LUT4 lut_inst_209 (
  .F(lut_f_209),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_209.INIT = 16'h8000;
LUT4 lut_inst_210 (
  .F(lut_f_210),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_210.INIT = 16'h8000;
LUT4 lut_inst_211 (
  .F(lut_f_211),
  .I0(lut_f_208),
  .I1(lut_f_209),
  .I2(lut_f_210),
  .I3(gw_vcc)
);
defparam lut_inst_211.INIT = 16'h8000;
LUT4 lut_inst_212 (
  .F(lut_f_212),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_212.INIT = 16'h8000;
LUT4 lut_inst_213 (
  .F(lut_f_213),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_213.INIT = 16'h8000;
LUT4 lut_inst_214 (
  .F(lut_f_214),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_214.INIT = 16'h8000;
LUT4 lut_inst_215 (
  .F(lut_f_215),
  .I0(lut_f_212),
  .I1(lut_f_213),
  .I2(lut_f_214),
  .I3(gw_vcc)
);
defparam lut_inst_215.INIT = 16'h8000;
LUT4 lut_inst_216 (
  .F(lut_f_216),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_216.INIT = 16'h8000;
LUT4 lut_inst_217 (
  .F(lut_f_217),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_217.INIT = 16'h8000;
LUT4 lut_inst_218 (
  .F(lut_f_218),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_218.INIT = 16'h8000;
LUT4 lut_inst_219 (
  .F(lut_f_219),
  .I0(lut_f_216),
  .I1(lut_f_217),
  .I2(lut_f_218),
  .I3(gw_vcc)
);
defparam lut_inst_219.INIT = 16'h8000;
LUT4 lut_inst_220 (
  .F(lut_f_220),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_220.INIT = 16'h8000;
LUT4 lut_inst_221 (
  .F(lut_f_221),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_221.INIT = 16'h8000;
LUT4 lut_inst_222 (
  .F(lut_f_222),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_222.INIT = 16'h8000;
LUT4 lut_inst_223 (
  .F(lut_f_223),
  .I0(lut_f_220),
  .I1(lut_f_221),
  .I2(lut_f_222),
  .I3(gw_vcc)
);
defparam lut_inst_223.INIT = 16'h8000;
LUT4 lut_inst_224 (
  .F(lut_f_224),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_224.INIT = 16'h8000;
LUT4 lut_inst_225 (
  .F(lut_f_225),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_225.INIT = 16'h8000;
LUT4 lut_inst_226 (
  .F(lut_f_226),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_226.INIT = 16'h8000;
LUT4 lut_inst_227 (
  .F(lut_f_227),
  .I0(lut_f_224),
  .I1(lut_f_225),
  .I2(lut_f_226),
  .I3(gw_vcc)
);
defparam lut_inst_227.INIT = 16'h8000;
LUT4 lut_inst_228 (
  .F(lut_f_228),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_228.INIT = 16'h8000;
LUT4 lut_inst_229 (
  .F(lut_f_229),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_229.INIT = 16'h8000;
LUT4 lut_inst_230 (
  .F(lut_f_230),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_230.INIT = 16'h8000;
LUT4 lut_inst_231 (
  .F(lut_f_231),
  .I0(lut_f_228),
  .I1(lut_f_229),
  .I2(lut_f_230),
  .I3(gw_vcc)
);
defparam lut_inst_231.INIT = 16'h8000;
LUT4 lut_inst_232 (
  .F(lut_f_232),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_232.INIT = 16'h8000;
LUT4 lut_inst_233 (
  .F(lut_f_233),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_233.INIT = 16'h8000;
LUT4 lut_inst_234 (
  .F(lut_f_234),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_234.INIT = 16'h8000;
LUT4 lut_inst_235 (
  .F(lut_f_235),
  .I0(lut_f_232),
  .I1(lut_f_233),
  .I2(lut_f_234),
  .I3(gw_vcc)
);
defparam lut_inst_235.INIT = 16'h8000;
LUT4 lut_inst_236 (
  .F(lut_f_236),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_236.INIT = 16'h8000;
LUT4 lut_inst_237 (
  .F(lut_f_237),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_237.INIT = 16'h8000;
LUT4 lut_inst_238 (
  .F(lut_f_238),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_238.INIT = 16'h8000;
LUT4 lut_inst_239 (
  .F(lut_f_239),
  .I0(lut_f_236),
  .I1(lut_f_237),
  .I2(lut_f_238),
  .I3(gw_vcc)
);
defparam lut_inst_239.INIT = 16'h8000;
LUT4 lut_inst_240 (
  .F(lut_f_240),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_240.INIT = 16'h8000;
LUT4 lut_inst_241 (
  .F(lut_f_241),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_241.INIT = 16'h8000;
LUT4 lut_inst_242 (
  .F(lut_f_242),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_242.INIT = 16'h8000;
LUT4 lut_inst_243 (
  .F(lut_f_243),
  .I0(lut_f_240),
  .I1(lut_f_241),
  .I2(lut_f_242),
  .I3(gw_vcc)
);
defparam lut_inst_243.INIT = 16'h8000;
LUT4 lut_inst_244 (
  .F(lut_f_244),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_244.INIT = 16'h8000;
LUT4 lut_inst_245 (
  .F(lut_f_245),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_245.INIT = 16'h8000;
LUT4 lut_inst_246 (
  .F(lut_f_246),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_246.INIT = 16'h8000;
LUT4 lut_inst_247 (
  .F(lut_f_247),
  .I0(lut_f_244),
  .I1(lut_f_245),
  .I2(lut_f_246),
  .I3(gw_vcc)
);
defparam lut_inst_247.INIT = 16'h8000;
LUT4 lut_inst_248 (
  .F(lut_f_248),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_248.INIT = 16'h8000;
LUT4 lut_inst_249 (
  .F(lut_f_249),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_249.INIT = 16'h8000;
LUT4 lut_inst_250 (
  .F(lut_f_250),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_250.INIT = 16'h8000;
LUT4 lut_inst_251 (
  .F(lut_f_251),
  .I0(lut_f_248),
  .I1(lut_f_249),
  .I2(lut_f_250),
  .I3(gw_vcc)
);
defparam lut_inst_251.INIT = 16'h8000;
LUT4 lut_inst_252 (
  .F(lut_f_252),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_252.INIT = 16'h8000;
LUT4 lut_inst_253 (
  .F(lut_f_253),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_253.INIT = 16'h8000;
LUT4 lut_inst_254 (
  .F(lut_f_254),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_254.INIT = 16'h8000;
LUT4 lut_inst_255 (
  .F(lut_f_255),
  .I0(lut_f_252),
  .I1(lut_f_253),
  .I2(lut_f_254),
  .I3(gw_vcc)
);
defparam lut_inst_255.INIT = 16'h8000;
LUT4 lut_inst_256 (
  .F(lut_f_256),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_256.INIT = 16'h8000;
LUT4 lut_inst_257 (
  .F(lut_f_257),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_257.INIT = 16'h8000;
LUT4 lut_inst_258 (
  .F(lut_f_258),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_258.INIT = 16'h8000;
LUT4 lut_inst_259 (
  .F(lut_f_259),
  .I0(lut_f_256),
  .I1(lut_f_257),
  .I2(lut_f_258),
  .I3(gw_vcc)
);
defparam lut_inst_259.INIT = 16'h8000;
LUT4 lut_inst_260 (
  .F(lut_f_260),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_260.INIT = 16'h8000;
LUT4 lut_inst_261 (
  .F(lut_f_261),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_261.INIT = 16'h8000;
LUT4 lut_inst_262 (
  .F(lut_f_262),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_262.INIT = 16'h8000;
LUT4 lut_inst_263 (
  .F(lut_f_263),
  .I0(lut_f_260),
  .I1(lut_f_261),
  .I2(lut_f_262),
  .I3(gw_vcc)
);
defparam lut_inst_263.INIT = 16'h8000;
LUT4 lut_inst_264 (
  .F(lut_f_264),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_264.INIT = 16'h8000;
LUT4 lut_inst_265 (
  .F(lut_f_265),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_265.INIT = 16'h8000;
LUT4 lut_inst_266 (
  .F(lut_f_266),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_266.INIT = 16'h8000;
LUT4 lut_inst_267 (
  .F(lut_f_267),
  .I0(lut_f_264),
  .I1(lut_f_265),
  .I2(lut_f_266),
  .I3(gw_vcc)
);
defparam lut_inst_267.INIT = 16'h8000;
LUT4 lut_inst_268 (
  .F(lut_f_268),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_268.INIT = 16'h8000;
LUT4 lut_inst_269 (
  .F(lut_f_269),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_269.INIT = 16'h8000;
LUT4 lut_inst_270 (
  .F(lut_f_270),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_270.INIT = 16'h8000;
LUT4 lut_inst_271 (
  .F(lut_f_271),
  .I0(lut_f_268),
  .I1(lut_f_269),
  .I2(lut_f_270),
  .I3(gw_vcc)
);
defparam lut_inst_271.INIT = 16'h8000;
LUT4 lut_inst_272 (
  .F(lut_f_272),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_272.INIT = 16'h8000;
LUT4 lut_inst_273 (
  .F(lut_f_273),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_273.INIT = 16'h8000;
LUT4 lut_inst_274 (
  .F(lut_f_274),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_274.INIT = 16'h8000;
LUT4 lut_inst_275 (
  .F(lut_f_275),
  .I0(lut_f_272),
  .I1(lut_f_273),
  .I2(lut_f_274),
  .I3(gw_vcc)
);
defparam lut_inst_275.INIT = 16'h8000;
LUT4 lut_inst_276 (
  .F(lut_f_276),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_276.INIT = 16'h8000;
LUT4 lut_inst_277 (
  .F(lut_f_277),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_277.INIT = 16'h8000;
LUT4 lut_inst_278 (
  .F(lut_f_278),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_278.INIT = 16'h8000;
LUT4 lut_inst_279 (
  .F(lut_f_279),
  .I0(lut_f_276),
  .I1(lut_f_277),
  .I2(lut_f_278),
  .I3(gw_vcc)
);
defparam lut_inst_279.INIT = 16'h8000;
LUT4 lut_inst_280 (
  .F(lut_f_280),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_280.INIT = 16'h8000;
LUT4 lut_inst_281 (
  .F(lut_f_281),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_281.INIT = 16'h8000;
LUT4 lut_inst_282 (
  .F(lut_f_282),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_282.INIT = 16'h8000;
LUT4 lut_inst_283 (
  .F(lut_f_283),
  .I0(lut_f_280),
  .I1(lut_f_281),
  .I2(lut_f_282),
  .I3(gw_vcc)
);
defparam lut_inst_283.INIT = 16'h8000;
LUT4 lut_inst_284 (
  .F(lut_f_284),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_284.INIT = 16'h8000;
LUT4 lut_inst_285 (
  .F(lut_f_285),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_285.INIT = 16'h8000;
LUT4 lut_inst_286 (
  .F(lut_f_286),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_286.INIT = 16'h8000;
LUT4 lut_inst_287 (
  .F(lut_f_287),
  .I0(lut_f_284),
  .I1(lut_f_285),
  .I2(lut_f_286),
  .I3(gw_vcc)
);
defparam lut_inst_287.INIT = 16'h8000;
LUT4 lut_inst_288 (
  .F(lut_f_288),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_288.INIT = 16'h8000;
LUT4 lut_inst_289 (
  .F(lut_f_289),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_289.INIT = 16'h8000;
LUT4 lut_inst_290 (
  .F(lut_f_290),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_290.INIT = 16'h8000;
LUT4 lut_inst_291 (
  .F(lut_f_291),
  .I0(lut_f_288),
  .I1(lut_f_289),
  .I2(lut_f_290),
  .I3(gw_vcc)
);
defparam lut_inst_291.INIT = 16'h8000;
LUT4 lut_inst_292 (
  .F(lut_f_292),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_292.INIT = 16'h8000;
LUT4 lut_inst_293 (
  .F(lut_f_293),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_293.INIT = 16'h8000;
LUT4 lut_inst_294 (
  .F(lut_f_294),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_294.INIT = 16'h8000;
LUT4 lut_inst_295 (
  .F(lut_f_295),
  .I0(lut_f_292),
  .I1(lut_f_293),
  .I2(lut_f_294),
  .I3(gw_vcc)
);
defparam lut_inst_295.INIT = 16'h8000;
LUT4 lut_inst_296 (
  .F(lut_f_296),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_296.INIT = 16'h8000;
LUT4 lut_inst_297 (
  .F(lut_f_297),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_297.INIT = 16'h8000;
LUT4 lut_inst_298 (
  .F(lut_f_298),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_298.INIT = 16'h8000;
LUT4 lut_inst_299 (
  .F(lut_f_299),
  .I0(lut_f_296),
  .I1(lut_f_297),
  .I2(lut_f_298),
  .I3(gw_vcc)
);
defparam lut_inst_299.INIT = 16'h8000;
LUT4 lut_inst_300 (
  .F(lut_f_300),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_300.INIT = 16'h8000;
LUT4 lut_inst_301 (
  .F(lut_f_301),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_301.INIT = 16'h8000;
LUT4 lut_inst_302 (
  .F(lut_f_302),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_302.INIT = 16'h8000;
LUT4 lut_inst_303 (
  .F(lut_f_303),
  .I0(lut_f_300),
  .I1(lut_f_301),
  .I2(lut_f_302),
  .I3(gw_vcc)
);
defparam lut_inst_303.INIT = 16'h8000;
LUT4 lut_inst_304 (
  .F(lut_f_304),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_304.INIT = 16'h8000;
LUT4 lut_inst_305 (
  .F(lut_f_305),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_305.INIT = 16'h8000;
LUT4 lut_inst_306 (
  .F(lut_f_306),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_306.INIT = 16'h8000;
LUT4 lut_inst_307 (
  .F(lut_f_307),
  .I0(lut_f_304),
  .I1(lut_f_305),
  .I2(lut_f_306),
  .I3(gw_vcc)
);
defparam lut_inst_307.INIT = 16'h8000;
LUT4 lut_inst_308 (
  .F(lut_f_308),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_308.INIT = 16'h8000;
LUT4 lut_inst_309 (
  .F(lut_f_309),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_309.INIT = 16'h8000;
LUT4 lut_inst_310 (
  .F(lut_f_310),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_310.INIT = 16'h8000;
LUT4 lut_inst_311 (
  .F(lut_f_311),
  .I0(lut_f_308),
  .I1(lut_f_309),
  .I2(lut_f_310),
  .I3(gw_vcc)
);
defparam lut_inst_311.INIT = 16'h8000;
LUT4 lut_inst_312 (
  .F(lut_f_312),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_312.INIT = 16'h8000;
LUT4 lut_inst_313 (
  .F(lut_f_313),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_313.INIT = 16'h8000;
LUT4 lut_inst_314 (
  .F(lut_f_314),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_314.INIT = 16'h8000;
LUT4 lut_inst_315 (
  .F(lut_f_315),
  .I0(lut_f_312),
  .I1(lut_f_313),
  .I2(lut_f_314),
  .I3(gw_vcc)
);
defparam lut_inst_315.INIT = 16'h8000;
LUT4 lut_inst_316 (
  .F(lut_f_316),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_316.INIT = 16'h8000;
LUT4 lut_inst_317 (
  .F(lut_f_317),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_317.INIT = 16'h8000;
LUT4 lut_inst_318 (
  .F(lut_f_318),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_318.INIT = 16'h8000;
LUT4 lut_inst_319 (
  .F(lut_f_319),
  .I0(lut_f_316),
  .I1(lut_f_317),
  .I2(lut_f_318),
  .I3(gw_vcc)
);
defparam lut_inst_319.INIT = 16'h8000;
LUT4 lut_inst_320 (
  .F(lut_f_320),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_320.INIT = 16'h8000;
LUT4 lut_inst_321 (
  .F(lut_f_321),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_321.INIT = 16'h8000;
LUT4 lut_inst_322 (
  .F(lut_f_322),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_322.INIT = 16'h8000;
LUT4 lut_inst_323 (
  .F(lut_f_323),
  .I0(lut_f_320),
  .I1(lut_f_321),
  .I2(lut_f_322),
  .I3(gw_vcc)
);
defparam lut_inst_323.INIT = 16'h8000;
LUT4 lut_inst_324 (
  .F(lut_f_324),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_324.INIT = 16'h8000;
LUT4 lut_inst_325 (
  .F(lut_f_325),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_325.INIT = 16'h8000;
LUT4 lut_inst_326 (
  .F(lut_f_326),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_326.INIT = 16'h8000;
LUT4 lut_inst_327 (
  .F(lut_f_327),
  .I0(lut_f_324),
  .I1(lut_f_325),
  .I2(lut_f_326),
  .I3(gw_vcc)
);
defparam lut_inst_327.INIT = 16'h8000;
LUT4 lut_inst_328 (
  .F(lut_f_328),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_328.INIT = 16'h8000;
LUT4 lut_inst_329 (
  .F(lut_f_329),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_329.INIT = 16'h8000;
LUT4 lut_inst_330 (
  .F(lut_f_330),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_330.INIT = 16'h8000;
LUT4 lut_inst_331 (
  .F(lut_f_331),
  .I0(lut_f_328),
  .I1(lut_f_329),
  .I2(lut_f_330),
  .I3(gw_vcc)
);
defparam lut_inst_331.INIT = 16'h8000;
LUT4 lut_inst_332 (
  .F(lut_f_332),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_332.INIT = 16'h8000;
LUT4 lut_inst_333 (
  .F(lut_f_333),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_333.INIT = 16'h8000;
LUT4 lut_inst_334 (
  .F(lut_f_334),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_334.INIT = 16'h8000;
LUT4 lut_inst_335 (
  .F(lut_f_335),
  .I0(lut_f_332),
  .I1(lut_f_333),
  .I2(lut_f_334),
  .I3(gw_vcc)
);
defparam lut_inst_335.INIT = 16'h8000;
LUT4 lut_inst_336 (
  .F(lut_f_336),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_336.INIT = 16'h8000;
LUT4 lut_inst_337 (
  .F(lut_f_337),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_337.INIT = 16'h8000;
LUT4 lut_inst_338 (
  .F(lut_f_338),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_338.INIT = 16'h8000;
LUT4 lut_inst_339 (
  .F(lut_f_339),
  .I0(lut_f_336),
  .I1(lut_f_337),
  .I2(lut_f_338),
  .I3(gw_vcc)
);
defparam lut_inst_339.INIT = 16'h8000;
LUT4 lut_inst_340 (
  .F(lut_f_340),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_340.INIT = 16'h8000;
LUT4 lut_inst_341 (
  .F(lut_f_341),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_341.INIT = 16'h8000;
LUT4 lut_inst_342 (
  .F(lut_f_342),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_342.INIT = 16'h8000;
LUT4 lut_inst_343 (
  .F(lut_f_343),
  .I0(lut_f_340),
  .I1(lut_f_341),
  .I2(lut_f_342),
  .I3(gw_vcc)
);
defparam lut_inst_343.INIT = 16'h8000;
LUT4 lut_inst_344 (
  .F(lut_f_344),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_344.INIT = 16'h8000;
LUT4 lut_inst_345 (
  .F(lut_f_345),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_345.INIT = 16'h8000;
LUT4 lut_inst_346 (
  .F(lut_f_346),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_346.INIT = 16'h8000;
LUT4 lut_inst_347 (
  .F(lut_f_347),
  .I0(lut_f_344),
  .I1(lut_f_345),
  .I2(lut_f_346),
  .I3(gw_vcc)
);
defparam lut_inst_347.INIT = 16'h8000;
LUT4 lut_inst_348 (
  .F(lut_f_348),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_348.INIT = 16'h8000;
LUT4 lut_inst_349 (
  .F(lut_f_349),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_349.INIT = 16'h8000;
LUT4 lut_inst_350 (
  .F(lut_f_350),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_350.INIT = 16'h8000;
LUT4 lut_inst_351 (
  .F(lut_f_351),
  .I0(lut_f_348),
  .I1(lut_f_349),
  .I2(lut_f_350),
  .I3(gw_vcc)
);
defparam lut_inst_351.INIT = 16'h8000;
LUT4 lut_inst_352 (
  .F(lut_f_352),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_352.INIT = 16'h8000;
LUT4 lut_inst_353 (
  .F(lut_f_353),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_353.INIT = 16'h8000;
LUT4 lut_inst_354 (
  .F(lut_f_354),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_354.INIT = 16'h8000;
LUT4 lut_inst_355 (
  .F(lut_f_355),
  .I0(lut_f_352),
  .I1(lut_f_353),
  .I2(lut_f_354),
  .I3(gw_vcc)
);
defparam lut_inst_355.INIT = 16'h8000;
LUT4 lut_inst_356 (
  .F(lut_f_356),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_356.INIT = 16'h8000;
LUT4 lut_inst_357 (
  .F(lut_f_357),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_357.INIT = 16'h8000;
LUT4 lut_inst_358 (
  .F(lut_f_358),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_358.INIT = 16'h8000;
LUT4 lut_inst_359 (
  .F(lut_f_359),
  .I0(lut_f_356),
  .I1(lut_f_357),
  .I2(lut_f_358),
  .I3(gw_vcc)
);
defparam lut_inst_359.INIT = 16'h8000;
LUT4 lut_inst_360 (
  .F(lut_f_360),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_360.INIT = 16'h8000;
LUT4 lut_inst_361 (
  .F(lut_f_361),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_361.INIT = 16'h8000;
LUT4 lut_inst_362 (
  .F(lut_f_362),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_362.INIT = 16'h8000;
LUT4 lut_inst_363 (
  .F(lut_f_363),
  .I0(lut_f_360),
  .I1(lut_f_361),
  .I2(lut_f_362),
  .I3(gw_vcc)
);
defparam lut_inst_363.INIT = 16'h8000;
LUT4 lut_inst_364 (
  .F(lut_f_364),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_364.INIT = 16'h8000;
LUT4 lut_inst_365 (
  .F(lut_f_365),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_365.INIT = 16'h8000;
LUT4 lut_inst_366 (
  .F(lut_f_366),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_366.INIT = 16'h8000;
LUT4 lut_inst_367 (
  .F(lut_f_367),
  .I0(lut_f_364),
  .I1(lut_f_365),
  .I2(lut_f_366),
  .I3(gw_vcc)
);
defparam lut_inst_367.INIT = 16'h8000;
LUT4 lut_inst_368 (
  .F(lut_f_368),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_368.INIT = 16'h8000;
LUT4 lut_inst_369 (
  .F(lut_f_369),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_369.INIT = 16'h8000;
LUT4 lut_inst_370 (
  .F(lut_f_370),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_370.INIT = 16'h8000;
LUT4 lut_inst_371 (
  .F(lut_f_371),
  .I0(lut_f_368),
  .I1(lut_f_369),
  .I2(lut_f_370),
  .I3(gw_vcc)
);
defparam lut_inst_371.INIT = 16'h8000;
LUT4 lut_inst_372 (
  .F(lut_f_372),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_372.INIT = 16'h8000;
LUT4 lut_inst_373 (
  .F(lut_f_373),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_373.INIT = 16'h8000;
LUT4 lut_inst_374 (
  .F(lut_f_374),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_374.INIT = 16'h8000;
LUT4 lut_inst_375 (
  .F(lut_f_375),
  .I0(lut_f_372),
  .I1(lut_f_373),
  .I2(lut_f_374),
  .I3(gw_vcc)
);
defparam lut_inst_375.INIT = 16'h8000;
LUT4 lut_inst_376 (
  .F(lut_f_376),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_376.INIT = 16'h8000;
LUT4 lut_inst_377 (
  .F(lut_f_377),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_377.INIT = 16'h8000;
LUT4 lut_inst_378 (
  .F(lut_f_378),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_378.INIT = 16'h8000;
LUT4 lut_inst_379 (
  .F(lut_f_379),
  .I0(lut_f_376),
  .I1(lut_f_377),
  .I2(lut_f_378),
  .I3(gw_vcc)
);
defparam lut_inst_379.INIT = 16'h8000;
LUT4 lut_inst_380 (
  .F(lut_f_380),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_380.INIT = 16'h8000;
LUT4 lut_inst_381 (
  .F(lut_f_381),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_381.INIT = 16'h8000;
LUT4 lut_inst_382 (
  .F(lut_f_382),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_382.INIT = 16'h8000;
LUT4 lut_inst_383 (
  .F(lut_f_383),
  .I0(lut_f_380),
  .I1(lut_f_381),
  .I2(lut_f_382),
  .I3(gw_vcc)
);
defparam lut_inst_383.INIT = 16'h8000;
LUT4 lut_inst_384 (
  .F(lut_f_384),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_384.INIT = 16'h8000;
LUT4 lut_inst_385 (
  .F(lut_f_385),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_385.INIT = 16'h8000;
LUT4 lut_inst_386 (
  .F(lut_f_386),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_386.INIT = 16'h8000;
LUT4 lut_inst_387 (
  .F(lut_f_387),
  .I0(lut_f_384),
  .I1(lut_f_385),
  .I2(lut_f_386),
  .I3(gw_vcc)
);
defparam lut_inst_387.INIT = 16'h8000;
LUT4 lut_inst_388 (
  .F(lut_f_388),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_388.INIT = 16'h8000;
LUT4 lut_inst_389 (
  .F(lut_f_389),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_389.INIT = 16'h8000;
LUT4 lut_inst_390 (
  .F(lut_f_390),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_390.INIT = 16'h8000;
LUT4 lut_inst_391 (
  .F(lut_f_391),
  .I0(lut_f_388),
  .I1(lut_f_389),
  .I2(lut_f_390),
  .I3(gw_vcc)
);
defparam lut_inst_391.INIT = 16'h8000;
LUT4 lut_inst_392 (
  .F(lut_f_392),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_392.INIT = 16'h8000;
LUT4 lut_inst_393 (
  .F(lut_f_393),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_393.INIT = 16'h8000;
LUT4 lut_inst_394 (
  .F(lut_f_394),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_394.INIT = 16'h8000;
LUT4 lut_inst_395 (
  .F(lut_f_395),
  .I0(lut_f_392),
  .I1(lut_f_393),
  .I2(lut_f_394),
  .I3(gw_vcc)
);
defparam lut_inst_395.INIT = 16'h8000;
LUT4 lut_inst_396 (
  .F(lut_f_396),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_396.INIT = 16'h8000;
LUT4 lut_inst_397 (
  .F(lut_f_397),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_397.INIT = 16'h8000;
LUT4 lut_inst_398 (
  .F(lut_f_398),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_398.INIT = 16'h8000;
LUT4 lut_inst_399 (
  .F(lut_f_399),
  .I0(lut_f_396),
  .I1(lut_f_397),
  .I2(lut_f_398),
  .I3(gw_vcc)
);
defparam lut_inst_399.INIT = 16'h8000;
LUT4 lut_inst_400 (
  .F(lut_f_400),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_400.INIT = 16'h8000;
LUT4 lut_inst_401 (
  .F(lut_f_401),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_401.INIT = 16'h8000;
LUT4 lut_inst_402 (
  .F(lut_f_402),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_402.INIT = 16'h8000;
LUT4 lut_inst_403 (
  .F(lut_f_403),
  .I0(lut_f_400),
  .I1(lut_f_401),
  .I2(lut_f_402),
  .I3(gw_vcc)
);
defparam lut_inst_403.INIT = 16'h8000;
LUT4 lut_inst_404 (
  .F(lut_f_404),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_404.INIT = 16'h8000;
LUT4 lut_inst_405 (
  .F(lut_f_405),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_405.INIT = 16'h8000;
LUT4 lut_inst_406 (
  .F(lut_f_406),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_406.INIT = 16'h8000;
LUT4 lut_inst_407 (
  .F(lut_f_407),
  .I0(lut_f_404),
  .I1(lut_f_405),
  .I2(lut_f_406),
  .I3(gw_vcc)
);
defparam lut_inst_407.INIT = 16'h8000;
LUT4 lut_inst_408 (
  .F(lut_f_408),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_408.INIT = 16'h8000;
LUT4 lut_inst_409 (
  .F(lut_f_409),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_409.INIT = 16'h8000;
LUT4 lut_inst_410 (
  .F(lut_f_410),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_410.INIT = 16'h8000;
LUT4 lut_inst_411 (
  .F(lut_f_411),
  .I0(lut_f_408),
  .I1(lut_f_409),
  .I2(lut_f_410),
  .I3(gw_vcc)
);
defparam lut_inst_411.INIT = 16'h8000;
LUT4 lut_inst_412 (
  .F(lut_f_412),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_412.INIT = 16'h8000;
LUT4 lut_inst_413 (
  .F(lut_f_413),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_413.INIT = 16'h8000;
LUT4 lut_inst_414 (
  .F(lut_f_414),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_414.INIT = 16'h8000;
LUT4 lut_inst_415 (
  .F(lut_f_415),
  .I0(lut_f_412),
  .I1(lut_f_413),
  .I2(lut_f_414),
  .I3(gw_vcc)
);
defparam lut_inst_415.INIT = 16'h8000;
LUT4 lut_inst_416 (
  .F(lut_f_416),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_416.INIT = 16'h8000;
LUT4 lut_inst_417 (
  .F(lut_f_417),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_417.INIT = 16'h8000;
LUT4 lut_inst_418 (
  .F(lut_f_418),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_418.INIT = 16'h8000;
LUT4 lut_inst_419 (
  .F(lut_f_419),
  .I0(lut_f_416),
  .I1(lut_f_417),
  .I2(lut_f_418),
  .I3(gw_vcc)
);
defparam lut_inst_419.INIT = 16'h8000;
LUT4 lut_inst_420 (
  .F(lut_f_420),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_420.INIT = 16'h8000;
LUT4 lut_inst_421 (
  .F(lut_f_421),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_421.INIT = 16'h8000;
LUT4 lut_inst_422 (
  .F(lut_f_422),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_422.INIT = 16'h8000;
LUT4 lut_inst_423 (
  .F(lut_f_423),
  .I0(lut_f_420),
  .I1(lut_f_421),
  .I2(lut_f_422),
  .I3(gw_vcc)
);
defparam lut_inst_423.INIT = 16'h8000;
LUT4 lut_inst_424 (
  .F(lut_f_424),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_424.INIT = 16'h8000;
LUT4 lut_inst_425 (
  .F(lut_f_425),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_425.INIT = 16'h8000;
LUT4 lut_inst_426 (
  .F(lut_f_426),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_426.INIT = 16'h8000;
LUT4 lut_inst_427 (
  .F(lut_f_427),
  .I0(lut_f_424),
  .I1(lut_f_425),
  .I2(lut_f_426),
  .I3(gw_vcc)
);
defparam lut_inst_427.INIT = 16'h8000;
LUT4 lut_inst_428 (
  .F(lut_f_428),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_428.INIT = 16'h8000;
LUT4 lut_inst_429 (
  .F(lut_f_429),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_429.INIT = 16'h8000;
LUT4 lut_inst_430 (
  .F(lut_f_430),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_430.INIT = 16'h8000;
LUT4 lut_inst_431 (
  .F(lut_f_431),
  .I0(lut_f_428),
  .I1(lut_f_429),
  .I2(lut_f_430),
  .I3(gw_vcc)
);
defparam lut_inst_431.INIT = 16'h8000;
LUT4 lut_inst_432 (
  .F(lut_f_432),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_432.INIT = 16'h8000;
LUT4 lut_inst_433 (
  .F(lut_f_433),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_433.INIT = 16'h8000;
LUT4 lut_inst_434 (
  .F(lut_f_434),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_434.INIT = 16'h8000;
LUT4 lut_inst_435 (
  .F(lut_f_435),
  .I0(lut_f_432),
  .I1(lut_f_433),
  .I2(lut_f_434),
  .I3(gw_vcc)
);
defparam lut_inst_435.INIT = 16'h8000;
LUT4 lut_inst_436 (
  .F(lut_f_436),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_436.INIT = 16'h8000;
LUT4 lut_inst_437 (
  .F(lut_f_437),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_437.INIT = 16'h8000;
LUT4 lut_inst_438 (
  .F(lut_f_438),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_438.INIT = 16'h8000;
LUT4 lut_inst_439 (
  .F(lut_f_439),
  .I0(lut_f_436),
  .I1(lut_f_437),
  .I2(lut_f_438),
  .I3(gw_vcc)
);
defparam lut_inst_439.INIT = 16'h8000;
LUT4 lut_inst_440 (
  .F(lut_f_440),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_440.INIT = 16'h8000;
LUT4 lut_inst_441 (
  .F(lut_f_441),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_441.INIT = 16'h8000;
LUT4 lut_inst_442 (
  .F(lut_f_442),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_442.INIT = 16'h8000;
LUT4 lut_inst_443 (
  .F(lut_f_443),
  .I0(lut_f_440),
  .I1(lut_f_441),
  .I2(lut_f_442),
  .I3(gw_vcc)
);
defparam lut_inst_443.INIT = 16'h8000;
LUT4 lut_inst_444 (
  .F(lut_f_444),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_444.INIT = 16'h8000;
LUT4 lut_inst_445 (
  .F(lut_f_445),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_445.INIT = 16'h8000;
LUT4 lut_inst_446 (
  .F(lut_f_446),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_446.INIT = 16'h8000;
LUT4 lut_inst_447 (
  .F(lut_f_447),
  .I0(lut_f_444),
  .I1(lut_f_445),
  .I2(lut_f_446),
  .I3(gw_vcc)
);
defparam lut_inst_447.INIT = 16'h8000;
LUT4 lut_inst_448 (
  .F(lut_f_448),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_448.INIT = 16'h8000;
LUT4 lut_inst_449 (
  .F(lut_f_449),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_449.INIT = 16'h8000;
LUT4 lut_inst_450 (
  .F(lut_f_450),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_450.INIT = 16'h8000;
LUT4 lut_inst_451 (
  .F(lut_f_451),
  .I0(lut_f_448),
  .I1(lut_f_449),
  .I2(lut_f_450),
  .I3(gw_vcc)
);
defparam lut_inst_451.INIT = 16'h8000;
LUT4 lut_inst_452 (
  .F(lut_f_452),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_452.INIT = 16'h8000;
LUT4 lut_inst_453 (
  .F(lut_f_453),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_453.INIT = 16'h8000;
LUT4 lut_inst_454 (
  .F(lut_f_454),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_454.INIT = 16'h8000;
LUT4 lut_inst_455 (
  .F(lut_f_455),
  .I0(lut_f_452),
  .I1(lut_f_453),
  .I2(lut_f_454),
  .I3(gw_vcc)
);
defparam lut_inst_455.INIT = 16'h8000;
LUT4 lut_inst_456 (
  .F(lut_f_456),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_456.INIT = 16'h8000;
LUT4 lut_inst_457 (
  .F(lut_f_457),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_457.INIT = 16'h8000;
LUT4 lut_inst_458 (
  .F(lut_f_458),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_458.INIT = 16'h8000;
LUT4 lut_inst_459 (
  .F(lut_f_459),
  .I0(lut_f_456),
  .I1(lut_f_457),
  .I2(lut_f_458),
  .I3(gw_vcc)
);
defparam lut_inst_459.INIT = 16'h8000;
LUT4 lut_inst_460 (
  .F(lut_f_460),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_460.INIT = 16'h8000;
LUT4 lut_inst_461 (
  .F(lut_f_461),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_461.INIT = 16'h8000;
LUT4 lut_inst_462 (
  .F(lut_f_462),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_462.INIT = 16'h8000;
LUT4 lut_inst_463 (
  .F(lut_f_463),
  .I0(lut_f_460),
  .I1(lut_f_461),
  .I2(lut_f_462),
  .I3(gw_vcc)
);
defparam lut_inst_463.INIT = 16'h8000;
LUT4 lut_inst_464 (
  .F(lut_f_464),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_464.INIT = 16'h8000;
LUT4 lut_inst_465 (
  .F(lut_f_465),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_465.INIT = 16'h8000;
LUT4 lut_inst_466 (
  .F(lut_f_466),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_466.INIT = 16'h8000;
LUT4 lut_inst_467 (
  .F(lut_f_467),
  .I0(lut_f_464),
  .I1(lut_f_465),
  .I2(lut_f_466),
  .I3(gw_vcc)
);
defparam lut_inst_467.INIT = 16'h8000;
LUT4 lut_inst_468 (
  .F(lut_f_468),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_468.INIT = 16'h8000;
LUT4 lut_inst_469 (
  .F(lut_f_469),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_469.INIT = 16'h8000;
LUT4 lut_inst_470 (
  .F(lut_f_470),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_470.INIT = 16'h8000;
LUT4 lut_inst_471 (
  .F(lut_f_471),
  .I0(lut_f_468),
  .I1(lut_f_469),
  .I2(lut_f_470),
  .I3(gw_vcc)
);
defparam lut_inst_471.INIT = 16'h8000;
LUT4 lut_inst_472 (
  .F(lut_f_472),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_472.INIT = 16'h8000;
LUT4 lut_inst_473 (
  .F(lut_f_473),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_473.INIT = 16'h8000;
LUT4 lut_inst_474 (
  .F(lut_f_474),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_474.INIT = 16'h8000;
LUT4 lut_inst_475 (
  .F(lut_f_475),
  .I0(lut_f_472),
  .I1(lut_f_473),
  .I2(lut_f_474),
  .I3(gw_vcc)
);
defparam lut_inst_475.INIT = 16'h8000;
LUT4 lut_inst_476 (
  .F(lut_f_476),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_476.INIT = 16'h8000;
LUT4 lut_inst_477 (
  .F(lut_f_477),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_477.INIT = 16'h8000;
LUT4 lut_inst_478 (
  .F(lut_f_478),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_478.INIT = 16'h8000;
LUT4 lut_inst_479 (
  .F(lut_f_479),
  .I0(lut_f_476),
  .I1(lut_f_477),
  .I2(lut_f_478),
  .I3(gw_vcc)
);
defparam lut_inst_479.INIT = 16'h8000;
LUT4 lut_inst_480 (
  .F(lut_f_480),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_480.INIT = 16'h8000;
LUT4 lut_inst_481 (
  .F(lut_f_481),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_481.INIT = 16'h8000;
LUT4 lut_inst_482 (
  .F(lut_f_482),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_482.INIT = 16'h8000;
LUT4 lut_inst_483 (
  .F(lut_f_483),
  .I0(lut_f_480),
  .I1(lut_f_481),
  .I2(lut_f_482),
  .I3(gw_vcc)
);
defparam lut_inst_483.INIT = 16'h8000;
LUT4 lut_inst_484 (
  .F(lut_f_484),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_484.INIT = 16'h8000;
LUT4 lut_inst_485 (
  .F(lut_f_485),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_485.INIT = 16'h8000;
LUT4 lut_inst_486 (
  .F(lut_f_486),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_486.INIT = 16'h8000;
LUT4 lut_inst_487 (
  .F(lut_f_487),
  .I0(lut_f_484),
  .I1(lut_f_485),
  .I2(lut_f_486),
  .I3(gw_vcc)
);
defparam lut_inst_487.INIT = 16'h8000;
LUT4 lut_inst_488 (
  .F(lut_f_488),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_488.INIT = 16'h8000;
LUT4 lut_inst_489 (
  .F(lut_f_489),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_489.INIT = 16'h8000;
LUT4 lut_inst_490 (
  .F(lut_f_490),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_490.INIT = 16'h8000;
LUT4 lut_inst_491 (
  .F(lut_f_491),
  .I0(lut_f_488),
  .I1(lut_f_489),
  .I2(lut_f_490),
  .I3(gw_vcc)
);
defparam lut_inst_491.INIT = 16'h8000;
LUT4 lut_inst_492 (
  .F(lut_f_492),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_492.INIT = 16'h8000;
LUT4 lut_inst_493 (
  .F(lut_f_493),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_493.INIT = 16'h8000;
LUT4 lut_inst_494 (
  .F(lut_f_494),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_494.INIT = 16'h8000;
LUT4 lut_inst_495 (
  .F(lut_f_495),
  .I0(lut_f_492),
  .I1(lut_f_493),
  .I2(lut_f_494),
  .I3(gw_vcc)
);
defparam lut_inst_495.INIT = 16'h8000;
LUT4 lut_inst_496 (
  .F(lut_f_496),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_496.INIT = 16'h8000;
LUT4 lut_inst_497 (
  .F(lut_f_497),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_497.INIT = 16'h8000;
LUT4 lut_inst_498 (
  .F(lut_f_498),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_498.INIT = 16'h8000;
LUT4 lut_inst_499 (
  .F(lut_f_499),
  .I0(lut_f_496),
  .I1(lut_f_497),
  .I2(lut_f_498),
  .I3(gw_vcc)
);
defparam lut_inst_499.INIT = 16'h8000;
LUT4 lut_inst_500 (
  .F(lut_f_500),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_500.INIT = 16'h8000;
LUT4 lut_inst_501 (
  .F(lut_f_501),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_501.INIT = 16'h8000;
LUT4 lut_inst_502 (
  .F(lut_f_502),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_502.INIT = 16'h8000;
LUT4 lut_inst_503 (
  .F(lut_f_503),
  .I0(lut_f_500),
  .I1(lut_f_501),
  .I2(lut_f_502),
  .I3(gw_vcc)
);
defparam lut_inst_503.INIT = 16'h8000;
LUT4 lut_inst_504 (
  .F(lut_f_504),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_504.INIT = 16'h8000;
LUT4 lut_inst_505 (
  .F(lut_f_505),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_505.INIT = 16'h8000;
LUT4 lut_inst_506 (
  .F(lut_f_506),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_506.INIT = 16'h8000;
LUT4 lut_inst_507 (
  .F(lut_f_507),
  .I0(lut_f_504),
  .I1(lut_f_505),
  .I2(lut_f_506),
  .I3(gw_vcc)
);
defparam lut_inst_507.INIT = 16'h8000;
LUT4 lut_inst_508 (
  .F(lut_f_508),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_508.INIT = 16'h8000;
LUT4 lut_inst_509 (
  .F(lut_f_509),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_509.INIT = 16'h8000;
LUT4 lut_inst_510 (
  .F(lut_f_510),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_510.INIT = 16'h8000;
LUT4 lut_inst_511 (
  .F(lut_f_511),
  .I0(lut_f_508),
  .I1(lut_f_509),
  .I2(lut_f_510),
  .I3(gw_vcc)
);
defparam lut_inst_511.INIT = 16'h8000;
LUT4 lut_inst_512 (
  .F(lut_f_512),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_512.INIT = 16'h8000;
LUT4 lut_inst_513 (
  .F(lut_f_513),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_513.INIT = 16'h8000;
LUT4 lut_inst_514 (
  .F(lut_f_514),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_514.INIT = 16'h8000;
LUT4 lut_inst_515 (
  .F(lut_f_515),
  .I0(lut_f_512),
  .I1(lut_f_513),
  .I2(lut_f_514),
  .I3(gw_vcc)
);
defparam lut_inst_515.INIT = 16'h8000;
LUT4 lut_inst_516 (
  .F(lut_f_516),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_516.INIT = 16'h8000;
LUT4 lut_inst_517 (
  .F(lut_f_517),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_517.INIT = 16'h8000;
LUT4 lut_inst_518 (
  .F(lut_f_518),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_518.INIT = 16'h8000;
LUT4 lut_inst_519 (
  .F(lut_f_519),
  .I0(lut_f_516),
  .I1(lut_f_517),
  .I2(lut_f_518),
  .I3(gw_vcc)
);
defparam lut_inst_519.INIT = 16'h8000;
LUT4 lut_inst_520 (
  .F(lut_f_520),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_520.INIT = 16'h8000;
LUT4 lut_inst_521 (
  .F(lut_f_521),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_521.INIT = 16'h8000;
LUT4 lut_inst_522 (
  .F(lut_f_522),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_522.INIT = 16'h8000;
LUT4 lut_inst_523 (
  .F(lut_f_523),
  .I0(lut_f_520),
  .I1(lut_f_521),
  .I2(lut_f_522),
  .I3(gw_vcc)
);
defparam lut_inst_523.INIT = 16'h8000;
LUT4 lut_inst_524 (
  .F(lut_f_524),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_524.INIT = 16'h8000;
LUT4 lut_inst_525 (
  .F(lut_f_525),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_525.INIT = 16'h8000;
LUT4 lut_inst_526 (
  .F(lut_f_526),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_526.INIT = 16'h8000;
LUT4 lut_inst_527 (
  .F(lut_f_527),
  .I0(lut_f_524),
  .I1(lut_f_525),
  .I2(lut_f_526),
  .I3(gw_vcc)
);
defparam lut_inst_527.INIT = 16'h8000;
LUT4 lut_inst_528 (
  .F(lut_f_528),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_528.INIT = 16'h8000;
LUT4 lut_inst_529 (
  .F(lut_f_529),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_529.INIT = 16'h8000;
LUT4 lut_inst_530 (
  .F(lut_f_530),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_530.INIT = 16'h8000;
LUT4 lut_inst_531 (
  .F(lut_f_531),
  .I0(lut_f_528),
  .I1(lut_f_529),
  .I2(lut_f_530),
  .I3(gw_vcc)
);
defparam lut_inst_531.INIT = 16'h8000;
LUT4 lut_inst_532 (
  .F(lut_f_532),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_532.INIT = 16'h8000;
LUT4 lut_inst_533 (
  .F(lut_f_533),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_533.INIT = 16'h8000;
LUT4 lut_inst_534 (
  .F(lut_f_534),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_534.INIT = 16'h8000;
LUT4 lut_inst_535 (
  .F(lut_f_535),
  .I0(lut_f_532),
  .I1(lut_f_533),
  .I2(lut_f_534),
  .I3(gw_vcc)
);
defparam lut_inst_535.INIT = 16'h8000;
LUT4 lut_inst_536 (
  .F(lut_f_536),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_536.INIT = 16'h8000;
LUT4 lut_inst_537 (
  .F(lut_f_537),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_537.INIT = 16'h8000;
LUT4 lut_inst_538 (
  .F(lut_f_538),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_538.INIT = 16'h8000;
LUT4 lut_inst_539 (
  .F(lut_f_539),
  .I0(lut_f_536),
  .I1(lut_f_537),
  .I2(lut_f_538),
  .I3(gw_vcc)
);
defparam lut_inst_539.INIT = 16'h8000;
LUT4 lut_inst_540 (
  .F(lut_f_540),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_540.INIT = 16'h8000;
LUT4 lut_inst_541 (
  .F(lut_f_541),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_541.INIT = 16'h8000;
LUT4 lut_inst_542 (
  .F(lut_f_542),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_542.INIT = 16'h8000;
LUT4 lut_inst_543 (
  .F(lut_f_543),
  .I0(lut_f_540),
  .I1(lut_f_541),
  .I2(lut_f_542),
  .I3(gw_vcc)
);
defparam lut_inst_543.INIT = 16'h8000;
LUT4 lut_inst_544 (
  .F(lut_f_544),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_544.INIT = 16'h8000;
LUT4 lut_inst_545 (
  .F(lut_f_545),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_545.INIT = 16'h8000;
LUT4 lut_inst_546 (
  .F(lut_f_546),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_546.INIT = 16'h8000;
LUT4 lut_inst_547 (
  .F(lut_f_547),
  .I0(lut_f_544),
  .I1(lut_f_545),
  .I2(lut_f_546),
  .I3(gw_vcc)
);
defparam lut_inst_547.INIT = 16'h8000;
LUT4 lut_inst_548 (
  .F(lut_f_548),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_548.INIT = 16'h8000;
LUT4 lut_inst_549 (
  .F(lut_f_549),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_549.INIT = 16'h8000;
LUT4 lut_inst_550 (
  .F(lut_f_550),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_550.INIT = 16'h8000;
LUT4 lut_inst_551 (
  .F(lut_f_551),
  .I0(lut_f_548),
  .I1(lut_f_549),
  .I2(lut_f_550),
  .I3(gw_vcc)
);
defparam lut_inst_551.INIT = 16'h8000;
LUT4 lut_inst_552 (
  .F(lut_f_552),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_552.INIT = 16'h8000;
LUT4 lut_inst_553 (
  .F(lut_f_553),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_553.INIT = 16'h8000;
LUT4 lut_inst_554 (
  .F(lut_f_554),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_554.INIT = 16'h8000;
LUT4 lut_inst_555 (
  .F(lut_f_555),
  .I0(lut_f_552),
  .I1(lut_f_553),
  .I2(lut_f_554),
  .I3(gw_vcc)
);
defparam lut_inst_555.INIT = 16'h8000;
LUT4 lut_inst_556 (
  .F(lut_f_556),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_556.INIT = 16'h8000;
LUT4 lut_inst_557 (
  .F(lut_f_557),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_557.INIT = 16'h8000;
LUT4 lut_inst_558 (
  .F(lut_f_558),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_558.INIT = 16'h8000;
LUT4 lut_inst_559 (
  .F(lut_f_559),
  .I0(lut_f_556),
  .I1(lut_f_557),
  .I2(lut_f_558),
  .I3(gw_vcc)
);
defparam lut_inst_559.INIT = 16'h8000;
LUT4 lut_inst_560 (
  .F(lut_f_560),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_560.INIT = 16'h8000;
LUT4 lut_inst_561 (
  .F(lut_f_561),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_561.INIT = 16'h8000;
LUT4 lut_inst_562 (
  .F(lut_f_562),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_562.INIT = 16'h8000;
LUT4 lut_inst_563 (
  .F(lut_f_563),
  .I0(lut_f_560),
  .I1(lut_f_561),
  .I2(lut_f_562),
  .I3(gw_vcc)
);
defparam lut_inst_563.INIT = 16'h8000;
LUT4 lut_inst_564 (
  .F(lut_f_564),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_564.INIT = 16'h8000;
LUT4 lut_inst_565 (
  .F(lut_f_565),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_565.INIT = 16'h8000;
LUT4 lut_inst_566 (
  .F(lut_f_566),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_566.INIT = 16'h8000;
LUT4 lut_inst_567 (
  .F(lut_f_567),
  .I0(lut_f_564),
  .I1(lut_f_565),
  .I2(lut_f_566),
  .I3(gw_vcc)
);
defparam lut_inst_567.INIT = 16'h8000;
LUT4 lut_inst_568 (
  .F(lut_f_568),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_568.INIT = 16'h8000;
LUT4 lut_inst_569 (
  .F(lut_f_569),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_569.INIT = 16'h8000;
LUT4 lut_inst_570 (
  .F(lut_f_570),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_570.INIT = 16'h8000;
LUT4 lut_inst_571 (
  .F(lut_f_571),
  .I0(lut_f_568),
  .I1(lut_f_569),
  .I2(lut_f_570),
  .I3(gw_vcc)
);
defparam lut_inst_571.INIT = 16'h8000;
LUT4 lut_inst_572 (
  .F(lut_f_572),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_572.INIT = 16'h8000;
LUT4 lut_inst_573 (
  .F(lut_f_573),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_573.INIT = 16'h8000;
LUT4 lut_inst_574 (
  .F(lut_f_574),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_574.INIT = 16'h8000;
LUT4 lut_inst_575 (
  .F(lut_f_575),
  .I0(lut_f_572),
  .I1(lut_f_573),
  .I2(lut_f_574),
  .I3(gw_vcc)
);
defparam lut_inst_575.INIT = 16'h8000;
LUT4 lut_inst_576 (
  .F(lut_f_576),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_576.INIT = 16'h8000;
LUT4 lut_inst_577 (
  .F(lut_f_577),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_577.INIT = 16'h8000;
LUT4 lut_inst_578 (
  .F(lut_f_578),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_578.INIT = 16'h8000;
LUT4 lut_inst_579 (
  .F(lut_f_579),
  .I0(lut_f_576),
  .I1(lut_f_577),
  .I2(lut_f_578),
  .I3(gw_vcc)
);
defparam lut_inst_579.INIT = 16'h8000;
LUT4 lut_inst_580 (
  .F(lut_f_580),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_580.INIT = 16'h8000;
LUT4 lut_inst_581 (
  .F(lut_f_581),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_581.INIT = 16'h8000;
LUT4 lut_inst_582 (
  .F(lut_f_582),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_582.INIT = 16'h8000;
LUT4 lut_inst_583 (
  .F(lut_f_583),
  .I0(lut_f_580),
  .I1(lut_f_581),
  .I2(lut_f_582),
  .I3(gw_vcc)
);
defparam lut_inst_583.INIT = 16'h8000;
LUT4 lut_inst_584 (
  .F(lut_f_584),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_584.INIT = 16'h8000;
LUT4 lut_inst_585 (
  .F(lut_f_585),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_585.INIT = 16'h8000;
LUT4 lut_inst_586 (
  .F(lut_f_586),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_586.INIT = 16'h8000;
LUT4 lut_inst_587 (
  .F(lut_f_587),
  .I0(lut_f_584),
  .I1(lut_f_585),
  .I2(lut_f_586),
  .I3(gw_vcc)
);
defparam lut_inst_587.INIT = 16'h8000;
LUT4 lut_inst_588 (
  .F(lut_f_588),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_588.INIT = 16'h8000;
LUT4 lut_inst_589 (
  .F(lut_f_589),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_589.INIT = 16'h8000;
LUT4 lut_inst_590 (
  .F(lut_f_590),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_590.INIT = 16'h8000;
LUT4 lut_inst_591 (
  .F(lut_f_591),
  .I0(lut_f_588),
  .I1(lut_f_589),
  .I2(lut_f_590),
  .I3(gw_vcc)
);
defparam lut_inst_591.INIT = 16'h8000;
LUT4 lut_inst_592 (
  .F(lut_f_592),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_592.INIT = 16'h8000;
LUT4 lut_inst_593 (
  .F(lut_f_593),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_593.INIT = 16'h8000;
LUT4 lut_inst_594 (
  .F(lut_f_594),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_594.INIT = 16'h8000;
LUT4 lut_inst_595 (
  .F(lut_f_595),
  .I0(lut_f_592),
  .I1(lut_f_593),
  .I2(lut_f_594),
  .I3(gw_vcc)
);
defparam lut_inst_595.INIT = 16'h8000;
LUT4 lut_inst_596 (
  .F(lut_f_596),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_596.INIT = 16'h8000;
LUT4 lut_inst_597 (
  .F(lut_f_597),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_597.INIT = 16'h8000;
LUT4 lut_inst_598 (
  .F(lut_f_598),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_598.INIT = 16'h8000;
LUT4 lut_inst_599 (
  .F(lut_f_599),
  .I0(lut_f_596),
  .I1(lut_f_597),
  .I2(lut_f_598),
  .I3(gw_vcc)
);
defparam lut_inst_599.INIT = 16'h8000;
LUT4 lut_inst_600 (
  .F(lut_f_600),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_600.INIT = 16'h8000;
LUT4 lut_inst_601 (
  .F(lut_f_601),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_601.INIT = 16'h8000;
LUT4 lut_inst_602 (
  .F(lut_f_602),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_602.INIT = 16'h8000;
LUT4 lut_inst_603 (
  .F(lut_f_603),
  .I0(lut_f_600),
  .I1(lut_f_601),
  .I2(lut_f_602),
  .I3(gw_vcc)
);
defparam lut_inst_603.INIT = 16'h8000;
LUT4 lut_inst_604 (
  .F(lut_f_604),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_604.INIT = 16'h8000;
LUT4 lut_inst_605 (
  .F(lut_f_605),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_605.INIT = 16'h8000;
LUT4 lut_inst_606 (
  .F(lut_f_606),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_606.INIT = 16'h8000;
LUT4 lut_inst_607 (
  .F(lut_f_607),
  .I0(lut_f_604),
  .I1(lut_f_605),
  .I2(lut_f_606),
  .I3(gw_vcc)
);
defparam lut_inst_607.INIT = 16'h8000;
LUT4 lut_inst_608 (
  .F(lut_f_608),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_608.INIT = 16'h8000;
LUT4 lut_inst_609 (
  .F(lut_f_609),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_609.INIT = 16'h8000;
LUT4 lut_inst_610 (
  .F(lut_f_610),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_610.INIT = 16'h8000;
LUT4 lut_inst_611 (
  .F(lut_f_611),
  .I0(lut_f_608),
  .I1(lut_f_609),
  .I2(lut_f_610),
  .I3(gw_vcc)
);
defparam lut_inst_611.INIT = 16'h8000;
LUT4 lut_inst_612 (
  .F(lut_f_612),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_612.INIT = 16'h8000;
LUT4 lut_inst_613 (
  .F(lut_f_613),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_613.INIT = 16'h8000;
LUT4 lut_inst_614 (
  .F(lut_f_614),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_614.INIT = 16'h8000;
LUT4 lut_inst_615 (
  .F(lut_f_615),
  .I0(lut_f_612),
  .I1(lut_f_613),
  .I2(lut_f_614),
  .I3(gw_vcc)
);
defparam lut_inst_615.INIT = 16'h8000;
LUT4 lut_inst_616 (
  .F(lut_f_616),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_616.INIT = 16'h8000;
LUT4 lut_inst_617 (
  .F(lut_f_617),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_617.INIT = 16'h8000;
LUT4 lut_inst_618 (
  .F(lut_f_618),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_618.INIT = 16'h8000;
LUT4 lut_inst_619 (
  .F(lut_f_619),
  .I0(lut_f_616),
  .I1(lut_f_617),
  .I2(lut_f_618),
  .I3(gw_vcc)
);
defparam lut_inst_619.INIT = 16'h8000;
LUT4 lut_inst_620 (
  .F(lut_f_620),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_620.INIT = 16'h8000;
LUT4 lut_inst_621 (
  .F(lut_f_621),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_621.INIT = 16'h8000;
LUT4 lut_inst_622 (
  .F(lut_f_622),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_622.INIT = 16'h8000;
LUT4 lut_inst_623 (
  .F(lut_f_623),
  .I0(lut_f_620),
  .I1(lut_f_621),
  .I2(lut_f_622),
  .I3(gw_vcc)
);
defparam lut_inst_623.INIT = 16'h8000;
LUT4 lut_inst_624 (
  .F(lut_f_624),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_624.INIT = 16'h8000;
LUT4 lut_inst_625 (
  .F(lut_f_625),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_625.INIT = 16'h8000;
LUT4 lut_inst_626 (
  .F(lut_f_626),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_626.INIT = 16'h8000;
LUT4 lut_inst_627 (
  .F(lut_f_627),
  .I0(lut_f_624),
  .I1(lut_f_625),
  .I2(lut_f_626),
  .I3(gw_vcc)
);
defparam lut_inst_627.INIT = 16'h8000;
LUT4 lut_inst_628 (
  .F(lut_f_628),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_628.INIT = 16'h8000;
LUT4 lut_inst_629 (
  .F(lut_f_629),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_629.INIT = 16'h8000;
LUT4 lut_inst_630 (
  .F(lut_f_630),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_630.INIT = 16'h8000;
LUT4 lut_inst_631 (
  .F(lut_f_631),
  .I0(lut_f_628),
  .I1(lut_f_629),
  .I2(lut_f_630),
  .I3(gw_vcc)
);
defparam lut_inst_631.INIT = 16'h8000;
LUT4 lut_inst_632 (
  .F(lut_f_632),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_632.INIT = 16'h8000;
LUT4 lut_inst_633 (
  .F(lut_f_633),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_633.INIT = 16'h8000;
LUT4 lut_inst_634 (
  .F(lut_f_634),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_634.INIT = 16'h8000;
LUT4 lut_inst_635 (
  .F(lut_f_635),
  .I0(lut_f_632),
  .I1(lut_f_633),
  .I2(lut_f_634),
  .I3(gw_vcc)
);
defparam lut_inst_635.INIT = 16'h8000;
LUT4 lut_inst_636 (
  .F(lut_f_636),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_636.INIT = 16'h8000;
LUT4 lut_inst_637 (
  .F(lut_f_637),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_637.INIT = 16'h8000;
LUT4 lut_inst_638 (
  .F(lut_f_638),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_638.INIT = 16'h8000;
LUT4 lut_inst_639 (
  .F(lut_f_639),
  .I0(lut_f_636),
  .I1(lut_f_637),
  .I2(lut_f_638),
  .I3(gw_vcc)
);
defparam lut_inst_639.INIT = 16'h8000;
LUT4 lut_inst_640 (
  .F(lut_f_640),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_640.INIT = 16'h8000;
LUT4 lut_inst_641 (
  .F(lut_f_641),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_641.INIT = 16'h8000;
LUT4 lut_inst_642 (
  .F(lut_f_642),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_642.INIT = 16'h8000;
LUT4 lut_inst_643 (
  .F(lut_f_643),
  .I0(lut_f_640),
  .I1(lut_f_641),
  .I2(lut_f_642),
  .I3(gw_vcc)
);
defparam lut_inst_643.INIT = 16'h8000;
LUT4 lut_inst_644 (
  .F(lut_f_644),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_644.INIT = 16'h8000;
LUT4 lut_inst_645 (
  .F(lut_f_645),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_645.INIT = 16'h8000;
LUT4 lut_inst_646 (
  .F(lut_f_646),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_646.INIT = 16'h8000;
LUT4 lut_inst_647 (
  .F(lut_f_647),
  .I0(lut_f_644),
  .I1(lut_f_645),
  .I2(lut_f_646),
  .I3(gw_vcc)
);
defparam lut_inst_647.INIT = 16'h8000;
LUT4 lut_inst_648 (
  .F(lut_f_648),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_648.INIT = 16'h8000;
LUT4 lut_inst_649 (
  .F(lut_f_649),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_649.INIT = 16'h8000;
LUT4 lut_inst_650 (
  .F(lut_f_650),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_650.INIT = 16'h8000;
LUT4 lut_inst_651 (
  .F(lut_f_651),
  .I0(lut_f_648),
  .I1(lut_f_649),
  .I2(lut_f_650),
  .I3(gw_vcc)
);
defparam lut_inst_651.INIT = 16'h8000;
LUT4 lut_inst_652 (
  .F(lut_f_652),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_652.INIT = 16'h8000;
LUT4 lut_inst_653 (
  .F(lut_f_653),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_653.INIT = 16'h8000;
LUT4 lut_inst_654 (
  .F(lut_f_654),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_654.INIT = 16'h8000;
LUT4 lut_inst_655 (
  .F(lut_f_655),
  .I0(lut_f_652),
  .I1(lut_f_653),
  .I2(lut_f_654),
  .I3(gw_vcc)
);
defparam lut_inst_655.INIT = 16'h8000;
LUT4 lut_inst_656 (
  .F(lut_f_656),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_656.INIT = 16'h8000;
LUT4 lut_inst_657 (
  .F(lut_f_657),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_657.INIT = 16'h8000;
LUT4 lut_inst_658 (
  .F(lut_f_658),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_658.INIT = 16'h8000;
LUT4 lut_inst_659 (
  .F(lut_f_659),
  .I0(lut_f_656),
  .I1(lut_f_657),
  .I2(lut_f_658),
  .I3(gw_vcc)
);
defparam lut_inst_659.INIT = 16'h8000;
LUT4 lut_inst_660 (
  .F(lut_f_660),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_660.INIT = 16'h8000;
LUT4 lut_inst_661 (
  .F(lut_f_661),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_661.INIT = 16'h8000;
LUT4 lut_inst_662 (
  .F(lut_f_662),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_662.INIT = 16'h8000;
LUT4 lut_inst_663 (
  .F(lut_f_663),
  .I0(lut_f_660),
  .I1(lut_f_661),
  .I2(lut_f_662),
  .I3(gw_vcc)
);
defparam lut_inst_663.INIT = 16'h8000;
LUT4 lut_inst_664 (
  .F(lut_f_664),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_664.INIT = 16'h8000;
LUT4 lut_inst_665 (
  .F(lut_f_665),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_665.INIT = 16'h8000;
LUT4 lut_inst_666 (
  .F(lut_f_666),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_666.INIT = 16'h8000;
LUT4 lut_inst_667 (
  .F(lut_f_667),
  .I0(lut_f_664),
  .I1(lut_f_665),
  .I2(lut_f_666),
  .I3(gw_vcc)
);
defparam lut_inst_667.INIT = 16'h8000;
LUT4 lut_inst_668 (
  .F(lut_f_668),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_668.INIT = 16'h8000;
LUT4 lut_inst_669 (
  .F(lut_f_669),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_669.INIT = 16'h8000;
LUT4 lut_inst_670 (
  .F(lut_f_670),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_670.INIT = 16'h8000;
LUT4 lut_inst_671 (
  .F(lut_f_671),
  .I0(lut_f_668),
  .I1(lut_f_669),
  .I2(lut_f_670),
  .I3(gw_vcc)
);
defparam lut_inst_671.INIT = 16'h8000;
LUT4 lut_inst_672 (
  .F(lut_f_672),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_672.INIT = 16'h8000;
LUT4 lut_inst_673 (
  .F(lut_f_673),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_673.INIT = 16'h8000;
LUT4 lut_inst_674 (
  .F(lut_f_674),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_674.INIT = 16'h8000;
LUT4 lut_inst_675 (
  .F(lut_f_675),
  .I0(lut_f_672),
  .I1(lut_f_673),
  .I2(lut_f_674),
  .I3(gw_vcc)
);
defparam lut_inst_675.INIT = 16'h8000;
LUT4 lut_inst_676 (
  .F(lut_f_676),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_676.INIT = 16'h8000;
LUT4 lut_inst_677 (
  .F(lut_f_677),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_677.INIT = 16'h8000;
LUT4 lut_inst_678 (
  .F(lut_f_678),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_678.INIT = 16'h8000;
LUT4 lut_inst_679 (
  .F(lut_f_679),
  .I0(lut_f_676),
  .I1(lut_f_677),
  .I2(lut_f_678),
  .I3(gw_vcc)
);
defparam lut_inst_679.INIT = 16'h8000;
LUT4 lut_inst_680 (
  .F(lut_f_680),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_680.INIT = 16'h8000;
LUT4 lut_inst_681 (
  .F(lut_f_681),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_681.INIT = 16'h8000;
LUT4 lut_inst_682 (
  .F(lut_f_682),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_682.INIT = 16'h8000;
LUT4 lut_inst_683 (
  .F(lut_f_683),
  .I0(lut_f_680),
  .I1(lut_f_681),
  .I2(lut_f_682),
  .I3(gw_vcc)
);
defparam lut_inst_683.INIT = 16'h8000;
LUT4 lut_inst_684 (
  .F(lut_f_684),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_684.INIT = 16'h8000;
LUT4 lut_inst_685 (
  .F(lut_f_685),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_685.INIT = 16'h8000;
LUT4 lut_inst_686 (
  .F(lut_f_686),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_686.INIT = 16'h8000;
LUT4 lut_inst_687 (
  .F(lut_f_687),
  .I0(lut_f_684),
  .I1(lut_f_685),
  .I2(lut_f_686),
  .I3(gw_vcc)
);
defparam lut_inst_687.INIT = 16'h8000;
LUT4 lut_inst_688 (
  .F(lut_f_688),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_688.INIT = 16'h8000;
LUT4 lut_inst_689 (
  .F(lut_f_689),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_689.INIT = 16'h8000;
LUT4 lut_inst_690 (
  .F(lut_f_690),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_690.INIT = 16'h8000;
LUT4 lut_inst_691 (
  .F(lut_f_691),
  .I0(lut_f_688),
  .I1(lut_f_689),
  .I2(lut_f_690),
  .I3(gw_vcc)
);
defparam lut_inst_691.INIT = 16'h8000;
LUT4 lut_inst_692 (
  .F(lut_f_692),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_692.INIT = 16'h8000;
LUT4 lut_inst_693 (
  .F(lut_f_693),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_693.INIT = 16'h8000;
LUT4 lut_inst_694 (
  .F(lut_f_694),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_694.INIT = 16'h8000;
LUT4 lut_inst_695 (
  .F(lut_f_695),
  .I0(lut_f_692),
  .I1(lut_f_693),
  .I2(lut_f_694),
  .I3(gw_vcc)
);
defparam lut_inst_695.INIT = 16'h8000;
LUT4 lut_inst_696 (
  .F(lut_f_696),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_696.INIT = 16'h8000;
LUT4 lut_inst_697 (
  .F(lut_f_697),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_697.INIT = 16'h8000;
LUT4 lut_inst_698 (
  .F(lut_f_698),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_698.INIT = 16'h8000;
LUT4 lut_inst_699 (
  .F(lut_f_699),
  .I0(lut_f_696),
  .I1(lut_f_697),
  .I2(lut_f_698),
  .I3(gw_vcc)
);
defparam lut_inst_699.INIT = 16'h8000;
LUT4 lut_inst_700 (
  .F(lut_f_700),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_700.INIT = 16'h8000;
LUT4 lut_inst_701 (
  .F(lut_f_701),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_701.INIT = 16'h8000;
LUT4 lut_inst_702 (
  .F(lut_f_702),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_702.INIT = 16'h8000;
LUT4 lut_inst_703 (
  .F(lut_f_703),
  .I0(lut_f_700),
  .I1(lut_f_701),
  .I2(lut_f_702),
  .I3(gw_vcc)
);
defparam lut_inst_703.INIT = 16'h8000;
LUT4 lut_inst_704 (
  .F(lut_f_704),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_704.INIT = 16'h8000;
LUT4 lut_inst_705 (
  .F(lut_f_705),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_705.INIT = 16'h8000;
LUT4 lut_inst_706 (
  .F(lut_f_706),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_706.INIT = 16'h8000;
LUT4 lut_inst_707 (
  .F(lut_f_707),
  .I0(lut_f_704),
  .I1(lut_f_705),
  .I2(lut_f_706),
  .I3(gw_vcc)
);
defparam lut_inst_707.INIT = 16'h8000;
LUT4 lut_inst_708 (
  .F(lut_f_708),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_708.INIT = 16'h8000;
LUT4 lut_inst_709 (
  .F(lut_f_709),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_709.INIT = 16'h8000;
LUT4 lut_inst_710 (
  .F(lut_f_710),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_710.INIT = 16'h8000;
LUT4 lut_inst_711 (
  .F(lut_f_711),
  .I0(lut_f_708),
  .I1(lut_f_709),
  .I2(lut_f_710),
  .I3(gw_vcc)
);
defparam lut_inst_711.INIT = 16'h8000;
LUT4 lut_inst_712 (
  .F(lut_f_712),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_712.INIT = 16'h8000;
LUT4 lut_inst_713 (
  .F(lut_f_713),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_713.INIT = 16'h8000;
LUT4 lut_inst_714 (
  .F(lut_f_714),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_714.INIT = 16'h8000;
LUT4 lut_inst_715 (
  .F(lut_f_715),
  .I0(lut_f_712),
  .I1(lut_f_713),
  .I2(lut_f_714),
  .I3(gw_vcc)
);
defparam lut_inst_715.INIT = 16'h8000;
LUT4 lut_inst_716 (
  .F(lut_f_716),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_716.INIT = 16'h8000;
LUT4 lut_inst_717 (
  .F(lut_f_717),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_717.INIT = 16'h8000;
LUT4 lut_inst_718 (
  .F(lut_f_718),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_718.INIT = 16'h8000;
LUT4 lut_inst_719 (
  .F(lut_f_719),
  .I0(lut_f_716),
  .I1(lut_f_717),
  .I2(lut_f_718),
  .I3(gw_vcc)
);
defparam lut_inst_719.INIT = 16'h8000;
LUT4 lut_inst_720 (
  .F(lut_f_720),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_720.INIT = 16'h8000;
LUT4 lut_inst_721 (
  .F(lut_f_721),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_721.INIT = 16'h8000;
LUT4 lut_inst_722 (
  .F(lut_f_722),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_722.INIT = 16'h8000;
LUT4 lut_inst_723 (
  .F(lut_f_723),
  .I0(lut_f_720),
  .I1(lut_f_721),
  .I2(lut_f_722),
  .I3(gw_vcc)
);
defparam lut_inst_723.INIT = 16'h8000;
LUT4 lut_inst_724 (
  .F(lut_f_724),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_724.INIT = 16'h8000;
LUT4 lut_inst_725 (
  .F(lut_f_725),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_725.INIT = 16'h8000;
LUT4 lut_inst_726 (
  .F(lut_f_726),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_726.INIT = 16'h8000;
LUT4 lut_inst_727 (
  .F(lut_f_727),
  .I0(lut_f_724),
  .I1(lut_f_725),
  .I2(lut_f_726),
  .I3(gw_vcc)
);
defparam lut_inst_727.INIT = 16'h8000;
LUT4 lut_inst_728 (
  .F(lut_f_728),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_728.INIT = 16'h8000;
LUT4 lut_inst_729 (
  .F(lut_f_729),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_729.INIT = 16'h8000;
LUT4 lut_inst_730 (
  .F(lut_f_730),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_730.INIT = 16'h8000;
LUT4 lut_inst_731 (
  .F(lut_f_731),
  .I0(lut_f_728),
  .I1(lut_f_729),
  .I2(lut_f_730),
  .I3(gw_vcc)
);
defparam lut_inst_731.INIT = 16'h8000;
LUT4 lut_inst_732 (
  .F(lut_f_732),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_732.INIT = 16'h8000;
LUT4 lut_inst_733 (
  .F(lut_f_733),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_733.INIT = 16'h8000;
LUT4 lut_inst_734 (
  .F(lut_f_734),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_734.INIT = 16'h8000;
LUT4 lut_inst_735 (
  .F(lut_f_735),
  .I0(lut_f_732),
  .I1(lut_f_733),
  .I2(lut_f_734),
  .I3(gw_vcc)
);
defparam lut_inst_735.INIT = 16'h8000;
LUT4 lut_inst_736 (
  .F(lut_f_736),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_736.INIT = 16'h8000;
LUT4 lut_inst_737 (
  .F(lut_f_737),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_737.INIT = 16'h8000;
LUT4 lut_inst_738 (
  .F(lut_f_738),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_738.INIT = 16'h8000;
LUT4 lut_inst_739 (
  .F(lut_f_739),
  .I0(lut_f_736),
  .I1(lut_f_737),
  .I2(lut_f_738),
  .I3(gw_vcc)
);
defparam lut_inst_739.INIT = 16'h8000;
LUT4 lut_inst_740 (
  .F(lut_f_740),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_740.INIT = 16'h8000;
LUT4 lut_inst_741 (
  .F(lut_f_741),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_741.INIT = 16'h8000;
LUT4 lut_inst_742 (
  .F(lut_f_742),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_742.INIT = 16'h8000;
LUT4 lut_inst_743 (
  .F(lut_f_743),
  .I0(lut_f_740),
  .I1(lut_f_741),
  .I2(lut_f_742),
  .I3(gw_vcc)
);
defparam lut_inst_743.INIT = 16'h8000;
LUT4 lut_inst_744 (
  .F(lut_f_744),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_744.INIT = 16'h8000;
LUT4 lut_inst_745 (
  .F(lut_f_745),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_745.INIT = 16'h8000;
LUT4 lut_inst_746 (
  .F(lut_f_746),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_746.INIT = 16'h8000;
LUT4 lut_inst_747 (
  .F(lut_f_747),
  .I0(lut_f_744),
  .I1(lut_f_745),
  .I2(lut_f_746),
  .I3(gw_vcc)
);
defparam lut_inst_747.INIT = 16'h8000;
LUT4 lut_inst_748 (
  .F(lut_f_748),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_748.INIT = 16'h8000;
LUT4 lut_inst_749 (
  .F(lut_f_749),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_749.INIT = 16'h8000;
LUT4 lut_inst_750 (
  .F(lut_f_750),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_750.INIT = 16'h8000;
LUT4 lut_inst_751 (
  .F(lut_f_751),
  .I0(lut_f_748),
  .I1(lut_f_749),
  .I2(lut_f_750),
  .I3(gw_vcc)
);
defparam lut_inst_751.INIT = 16'h8000;
LUT4 lut_inst_752 (
  .F(lut_f_752),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_752.INIT = 16'h8000;
LUT4 lut_inst_753 (
  .F(lut_f_753),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_753.INIT = 16'h8000;
LUT4 lut_inst_754 (
  .F(lut_f_754),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_754.INIT = 16'h8000;
LUT4 lut_inst_755 (
  .F(lut_f_755),
  .I0(lut_f_752),
  .I1(lut_f_753),
  .I2(lut_f_754),
  .I3(gw_vcc)
);
defparam lut_inst_755.INIT = 16'h8000;
LUT4 lut_inst_756 (
  .F(lut_f_756),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_756.INIT = 16'h8000;
LUT4 lut_inst_757 (
  .F(lut_f_757),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_757.INIT = 16'h8000;
LUT4 lut_inst_758 (
  .F(lut_f_758),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_758.INIT = 16'h8000;
LUT4 lut_inst_759 (
  .F(lut_f_759),
  .I0(lut_f_756),
  .I1(lut_f_757),
  .I2(lut_f_758),
  .I3(gw_vcc)
);
defparam lut_inst_759.INIT = 16'h8000;
LUT4 lut_inst_760 (
  .F(lut_f_760),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_760.INIT = 16'h8000;
LUT4 lut_inst_761 (
  .F(lut_f_761),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_761.INIT = 16'h8000;
LUT4 lut_inst_762 (
  .F(lut_f_762),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_762.INIT = 16'h8000;
LUT4 lut_inst_763 (
  .F(lut_f_763),
  .I0(lut_f_760),
  .I1(lut_f_761),
  .I2(lut_f_762),
  .I3(gw_vcc)
);
defparam lut_inst_763.INIT = 16'h8000;
LUT4 lut_inst_764 (
  .F(lut_f_764),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_764.INIT = 16'h8000;
LUT4 lut_inst_765 (
  .F(lut_f_765),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_765.INIT = 16'h8000;
LUT4 lut_inst_766 (
  .F(lut_f_766),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_766.INIT = 16'h8000;
LUT4 lut_inst_767 (
  .F(lut_f_767),
  .I0(lut_f_764),
  .I1(lut_f_765),
  .I2(lut_f_766),
  .I3(gw_vcc)
);
defparam lut_inst_767.INIT = 16'h8000;
LUT4 lut_inst_768 (
  .F(lut_f_768),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_768.INIT = 16'h8000;
LUT4 lut_inst_769 (
  .F(lut_f_769),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_769.INIT = 16'h8000;
LUT4 lut_inst_770 (
  .F(lut_f_770),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_770.INIT = 16'h8000;
LUT4 lut_inst_771 (
  .F(lut_f_771),
  .I0(lut_f_768),
  .I1(lut_f_769),
  .I2(lut_f_770),
  .I3(gw_vcc)
);
defparam lut_inst_771.INIT = 16'h8000;
LUT4 lut_inst_772 (
  .F(lut_f_772),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_772.INIT = 16'h8000;
LUT4 lut_inst_773 (
  .F(lut_f_773),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_773.INIT = 16'h8000;
LUT4 lut_inst_774 (
  .F(lut_f_774),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_774.INIT = 16'h8000;
LUT4 lut_inst_775 (
  .F(lut_f_775),
  .I0(lut_f_772),
  .I1(lut_f_773),
  .I2(lut_f_774),
  .I3(gw_vcc)
);
defparam lut_inst_775.INIT = 16'h8000;
LUT4 lut_inst_776 (
  .F(lut_f_776),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_776.INIT = 16'h8000;
LUT4 lut_inst_777 (
  .F(lut_f_777),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_777.INIT = 16'h8000;
LUT4 lut_inst_778 (
  .F(lut_f_778),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_778.INIT = 16'h8000;
LUT4 lut_inst_779 (
  .F(lut_f_779),
  .I0(lut_f_776),
  .I1(lut_f_777),
  .I2(lut_f_778),
  .I3(gw_vcc)
);
defparam lut_inst_779.INIT = 16'h8000;
LUT4 lut_inst_780 (
  .F(lut_f_780),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_780.INIT = 16'h8000;
LUT4 lut_inst_781 (
  .F(lut_f_781),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_781.INIT = 16'h8000;
LUT4 lut_inst_782 (
  .F(lut_f_782),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_782.INIT = 16'h8000;
LUT4 lut_inst_783 (
  .F(lut_f_783),
  .I0(lut_f_780),
  .I1(lut_f_781),
  .I2(lut_f_782),
  .I3(gw_vcc)
);
defparam lut_inst_783.INIT = 16'h8000;
LUT4 lut_inst_784 (
  .F(lut_f_784),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_784.INIT = 16'h8000;
LUT4 lut_inst_785 (
  .F(lut_f_785),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_785.INIT = 16'h8000;
LUT4 lut_inst_786 (
  .F(lut_f_786),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_786.INIT = 16'h8000;
LUT4 lut_inst_787 (
  .F(lut_f_787),
  .I0(lut_f_784),
  .I1(lut_f_785),
  .I2(lut_f_786),
  .I3(gw_vcc)
);
defparam lut_inst_787.INIT = 16'h8000;
LUT4 lut_inst_788 (
  .F(lut_f_788),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_788.INIT = 16'h8000;
LUT4 lut_inst_789 (
  .F(lut_f_789),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_789.INIT = 16'h8000;
LUT4 lut_inst_790 (
  .F(lut_f_790),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_790.INIT = 16'h8000;
LUT4 lut_inst_791 (
  .F(lut_f_791),
  .I0(lut_f_788),
  .I1(lut_f_789),
  .I2(lut_f_790),
  .I3(gw_vcc)
);
defparam lut_inst_791.INIT = 16'h8000;
LUT4 lut_inst_792 (
  .F(lut_f_792),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_792.INIT = 16'h8000;
LUT4 lut_inst_793 (
  .F(lut_f_793),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_793.INIT = 16'h8000;
LUT4 lut_inst_794 (
  .F(lut_f_794),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_794.INIT = 16'h8000;
LUT4 lut_inst_795 (
  .F(lut_f_795),
  .I0(lut_f_792),
  .I1(lut_f_793),
  .I2(lut_f_794),
  .I3(gw_vcc)
);
defparam lut_inst_795.INIT = 16'h8000;
LUT4 lut_inst_796 (
  .F(lut_f_796),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_796.INIT = 16'h8000;
LUT4 lut_inst_797 (
  .F(lut_f_797),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_797.INIT = 16'h8000;
LUT4 lut_inst_798 (
  .F(lut_f_798),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_798.INIT = 16'h8000;
LUT4 lut_inst_799 (
  .F(lut_f_799),
  .I0(lut_f_796),
  .I1(lut_f_797),
  .I2(lut_f_798),
  .I3(gw_vcc)
);
defparam lut_inst_799.INIT = 16'h8000;
LUT4 lut_inst_800 (
  .F(lut_f_800),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_800.INIT = 16'h8000;
LUT4 lut_inst_801 (
  .F(lut_f_801),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_801.INIT = 16'h8000;
LUT4 lut_inst_802 (
  .F(lut_f_802),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_802.INIT = 16'h8000;
LUT4 lut_inst_803 (
  .F(lut_f_803),
  .I0(lut_f_800),
  .I1(lut_f_801),
  .I2(lut_f_802),
  .I3(gw_vcc)
);
defparam lut_inst_803.INIT = 16'h8000;
LUT4 lut_inst_804 (
  .F(lut_f_804),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_804.INIT = 16'h8000;
LUT4 lut_inst_805 (
  .F(lut_f_805),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_805.INIT = 16'h8000;
LUT4 lut_inst_806 (
  .F(lut_f_806),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_806.INIT = 16'h8000;
LUT4 lut_inst_807 (
  .F(lut_f_807),
  .I0(lut_f_804),
  .I1(lut_f_805),
  .I2(lut_f_806),
  .I3(gw_vcc)
);
defparam lut_inst_807.INIT = 16'h8000;
LUT4 lut_inst_808 (
  .F(lut_f_808),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_808.INIT = 16'h8000;
LUT4 lut_inst_809 (
  .F(lut_f_809),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_809.INIT = 16'h8000;
LUT4 lut_inst_810 (
  .F(lut_f_810),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_810.INIT = 16'h8000;
LUT4 lut_inst_811 (
  .F(lut_f_811),
  .I0(lut_f_808),
  .I1(lut_f_809),
  .I2(lut_f_810),
  .I3(gw_vcc)
);
defparam lut_inst_811.INIT = 16'h8000;
LUT4 lut_inst_812 (
  .F(lut_f_812),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_812.INIT = 16'h8000;
LUT4 lut_inst_813 (
  .F(lut_f_813),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_813.INIT = 16'h8000;
LUT4 lut_inst_814 (
  .F(lut_f_814),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_814.INIT = 16'h8000;
LUT4 lut_inst_815 (
  .F(lut_f_815),
  .I0(lut_f_812),
  .I1(lut_f_813),
  .I2(lut_f_814),
  .I3(gw_vcc)
);
defparam lut_inst_815.INIT = 16'h8000;
LUT4 lut_inst_816 (
  .F(lut_f_816),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_816.INIT = 16'h8000;
LUT4 lut_inst_817 (
  .F(lut_f_817),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_817.INIT = 16'h8000;
LUT4 lut_inst_818 (
  .F(lut_f_818),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_818.INIT = 16'h8000;
LUT4 lut_inst_819 (
  .F(lut_f_819),
  .I0(lut_f_816),
  .I1(lut_f_817),
  .I2(lut_f_818),
  .I3(gw_vcc)
);
defparam lut_inst_819.INIT = 16'h8000;
LUT4 lut_inst_820 (
  .F(lut_f_820),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_820.INIT = 16'h8000;
LUT4 lut_inst_821 (
  .F(lut_f_821),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_821.INIT = 16'h8000;
LUT4 lut_inst_822 (
  .F(lut_f_822),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_822.INIT = 16'h8000;
LUT4 lut_inst_823 (
  .F(lut_f_823),
  .I0(lut_f_820),
  .I1(lut_f_821),
  .I2(lut_f_822),
  .I3(gw_vcc)
);
defparam lut_inst_823.INIT = 16'h8000;
LUT4 lut_inst_824 (
  .F(lut_f_824),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_824.INIT = 16'h8000;
LUT4 lut_inst_825 (
  .F(lut_f_825),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_825.INIT = 16'h8000;
LUT4 lut_inst_826 (
  .F(lut_f_826),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_826.INIT = 16'h8000;
LUT4 lut_inst_827 (
  .F(lut_f_827),
  .I0(lut_f_824),
  .I1(lut_f_825),
  .I2(lut_f_826),
  .I3(gw_vcc)
);
defparam lut_inst_827.INIT = 16'h8000;
LUT4 lut_inst_828 (
  .F(lut_f_828),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_828.INIT = 16'h8000;
LUT4 lut_inst_829 (
  .F(lut_f_829),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_829.INIT = 16'h8000;
LUT4 lut_inst_830 (
  .F(lut_f_830),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_830.INIT = 16'h8000;
LUT4 lut_inst_831 (
  .F(lut_f_831),
  .I0(lut_f_828),
  .I1(lut_f_829),
  .I2(lut_f_830),
  .I3(gw_vcc)
);
defparam lut_inst_831.INIT = 16'h8000;
LUT4 lut_inst_832 (
  .F(lut_f_832),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_832.INIT = 16'h8000;
LUT4 lut_inst_833 (
  .F(lut_f_833),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_833.INIT = 16'h8000;
LUT4 lut_inst_834 (
  .F(lut_f_834),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_834.INIT = 16'h8000;
LUT4 lut_inst_835 (
  .F(lut_f_835),
  .I0(lut_f_832),
  .I1(lut_f_833),
  .I2(lut_f_834),
  .I3(gw_vcc)
);
defparam lut_inst_835.INIT = 16'h8000;
LUT4 lut_inst_836 (
  .F(lut_f_836),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_836.INIT = 16'h8000;
LUT4 lut_inst_837 (
  .F(lut_f_837),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_837.INIT = 16'h8000;
LUT4 lut_inst_838 (
  .F(lut_f_838),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_838.INIT = 16'h8000;
LUT4 lut_inst_839 (
  .F(lut_f_839),
  .I0(lut_f_836),
  .I1(lut_f_837),
  .I2(lut_f_838),
  .I3(gw_vcc)
);
defparam lut_inst_839.INIT = 16'h8000;
LUT4 lut_inst_840 (
  .F(lut_f_840),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_840.INIT = 16'h8000;
LUT4 lut_inst_841 (
  .F(lut_f_841),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_841.INIT = 16'h8000;
LUT4 lut_inst_842 (
  .F(lut_f_842),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_842.INIT = 16'h8000;
LUT4 lut_inst_843 (
  .F(lut_f_843),
  .I0(lut_f_840),
  .I1(lut_f_841),
  .I2(lut_f_842),
  .I3(gw_vcc)
);
defparam lut_inst_843.INIT = 16'h8000;
LUT4 lut_inst_844 (
  .F(lut_f_844),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_844.INIT = 16'h8000;
LUT4 lut_inst_845 (
  .F(lut_f_845),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_845.INIT = 16'h8000;
LUT4 lut_inst_846 (
  .F(lut_f_846),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_846.INIT = 16'h8000;
LUT4 lut_inst_847 (
  .F(lut_f_847),
  .I0(lut_f_844),
  .I1(lut_f_845),
  .I2(lut_f_846),
  .I3(gw_vcc)
);
defparam lut_inst_847.INIT = 16'h8000;
LUT4 lut_inst_848 (
  .F(lut_f_848),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_848.INIT = 16'h8000;
LUT4 lut_inst_849 (
  .F(lut_f_849),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_849.INIT = 16'h8000;
LUT4 lut_inst_850 (
  .F(lut_f_850),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_850.INIT = 16'h8000;
LUT4 lut_inst_851 (
  .F(lut_f_851),
  .I0(lut_f_848),
  .I1(lut_f_849),
  .I2(lut_f_850),
  .I3(gw_vcc)
);
defparam lut_inst_851.INIT = 16'h8000;
LUT4 lut_inst_852 (
  .F(lut_f_852),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_852.INIT = 16'h8000;
LUT4 lut_inst_853 (
  .F(lut_f_853),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_853.INIT = 16'h8000;
LUT4 lut_inst_854 (
  .F(lut_f_854),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_854.INIT = 16'h8000;
LUT4 lut_inst_855 (
  .F(lut_f_855),
  .I0(lut_f_852),
  .I1(lut_f_853),
  .I2(lut_f_854),
  .I3(gw_vcc)
);
defparam lut_inst_855.INIT = 16'h8000;
LUT4 lut_inst_856 (
  .F(lut_f_856),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_856.INIT = 16'h8000;
LUT4 lut_inst_857 (
  .F(lut_f_857),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_857.INIT = 16'h8000;
LUT4 lut_inst_858 (
  .F(lut_f_858),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_858.INIT = 16'h8000;
LUT4 lut_inst_859 (
  .F(lut_f_859),
  .I0(lut_f_856),
  .I1(lut_f_857),
  .I2(lut_f_858),
  .I3(gw_vcc)
);
defparam lut_inst_859.INIT = 16'h8000;
LUT4 lut_inst_860 (
  .F(lut_f_860),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_860.INIT = 16'h8000;
LUT4 lut_inst_861 (
  .F(lut_f_861),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_861.INIT = 16'h8000;
LUT4 lut_inst_862 (
  .F(lut_f_862),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_862.INIT = 16'h8000;
LUT4 lut_inst_863 (
  .F(lut_f_863),
  .I0(lut_f_860),
  .I1(lut_f_861),
  .I2(lut_f_862),
  .I3(gw_vcc)
);
defparam lut_inst_863.INIT = 16'h8000;
LUT4 lut_inst_864 (
  .F(lut_f_864),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_864.INIT = 16'h8000;
LUT4 lut_inst_865 (
  .F(lut_f_865),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_865.INIT = 16'h8000;
LUT4 lut_inst_866 (
  .F(lut_f_866),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_866.INIT = 16'h8000;
LUT4 lut_inst_867 (
  .F(lut_f_867),
  .I0(lut_f_864),
  .I1(lut_f_865),
  .I2(lut_f_866),
  .I3(gw_vcc)
);
defparam lut_inst_867.INIT = 16'h8000;
LUT4 lut_inst_868 (
  .F(lut_f_868),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_868.INIT = 16'h8000;
LUT4 lut_inst_869 (
  .F(lut_f_869),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_869.INIT = 16'h8000;
LUT4 lut_inst_870 (
  .F(lut_f_870),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_870.INIT = 16'h8000;
LUT4 lut_inst_871 (
  .F(lut_f_871),
  .I0(lut_f_868),
  .I1(lut_f_869),
  .I2(lut_f_870),
  .I3(gw_vcc)
);
defparam lut_inst_871.INIT = 16'h8000;
LUT4 lut_inst_872 (
  .F(lut_f_872),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_872.INIT = 16'h8000;
LUT4 lut_inst_873 (
  .F(lut_f_873),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_873.INIT = 16'h8000;
LUT4 lut_inst_874 (
  .F(lut_f_874),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_874.INIT = 16'h8000;
LUT4 lut_inst_875 (
  .F(lut_f_875),
  .I0(lut_f_872),
  .I1(lut_f_873),
  .I2(lut_f_874),
  .I3(gw_vcc)
);
defparam lut_inst_875.INIT = 16'h8000;
LUT4 lut_inst_876 (
  .F(lut_f_876),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_876.INIT = 16'h8000;
LUT4 lut_inst_877 (
  .F(lut_f_877),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_877.INIT = 16'h8000;
LUT4 lut_inst_878 (
  .F(lut_f_878),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_878.INIT = 16'h8000;
LUT4 lut_inst_879 (
  .F(lut_f_879),
  .I0(lut_f_876),
  .I1(lut_f_877),
  .I2(lut_f_878),
  .I3(gw_vcc)
);
defparam lut_inst_879.INIT = 16'h8000;
LUT4 lut_inst_880 (
  .F(lut_f_880),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_880.INIT = 16'h8000;
LUT4 lut_inst_881 (
  .F(lut_f_881),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_881.INIT = 16'h8000;
LUT4 lut_inst_882 (
  .F(lut_f_882),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_882.INIT = 16'h8000;
LUT4 lut_inst_883 (
  .F(lut_f_883),
  .I0(lut_f_880),
  .I1(lut_f_881),
  .I2(lut_f_882),
  .I3(gw_vcc)
);
defparam lut_inst_883.INIT = 16'h8000;
LUT4 lut_inst_884 (
  .F(lut_f_884),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_884.INIT = 16'h8000;
LUT4 lut_inst_885 (
  .F(lut_f_885),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_885.INIT = 16'h8000;
LUT4 lut_inst_886 (
  .F(lut_f_886),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_886.INIT = 16'h8000;
LUT4 lut_inst_887 (
  .F(lut_f_887),
  .I0(lut_f_884),
  .I1(lut_f_885),
  .I2(lut_f_886),
  .I3(gw_vcc)
);
defparam lut_inst_887.INIT = 16'h8000;
LUT4 lut_inst_888 (
  .F(lut_f_888),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_888.INIT = 16'h8000;
LUT4 lut_inst_889 (
  .F(lut_f_889),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_889.INIT = 16'h8000;
LUT4 lut_inst_890 (
  .F(lut_f_890),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_890.INIT = 16'h8000;
LUT4 lut_inst_891 (
  .F(lut_f_891),
  .I0(lut_f_888),
  .I1(lut_f_889),
  .I2(lut_f_890),
  .I3(gw_vcc)
);
defparam lut_inst_891.INIT = 16'h8000;
LUT4 lut_inst_892 (
  .F(lut_f_892),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_892.INIT = 16'h8000;
LUT4 lut_inst_893 (
  .F(lut_f_893),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_893.INIT = 16'h8000;
LUT4 lut_inst_894 (
  .F(lut_f_894),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_894.INIT = 16'h8000;
LUT4 lut_inst_895 (
  .F(lut_f_895),
  .I0(lut_f_892),
  .I1(lut_f_893),
  .I2(lut_f_894),
  .I3(gw_vcc)
);
defparam lut_inst_895.INIT = 16'h8000;
LUT4 lut_inst_896 (
  .F(lut_f_896),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_896.INIT = 16'h8000;
LUT4 lut_inst_897 (
  .F(lut_f_897),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_897.INIT = 16'h8000;
LUT4 lut_inst_898 (
  .F(lut_f_898),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_898.INIT = 16'h8000;
LUT4 lut_inst_899 (
  .F(lut_f_899),
  .I0(lut_f_896),
  .I1(lut_f_897),
  .I2(lut_f_898),
  .I3(gw_vcc)
);
defparam lut_inst_899.INIT = 16'h8000;
LUT4 lut_inst_900 (
  .F(lut_f_900),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_900.INIT = 16'h8000;
LUT4 lut_inst_901 (
  .F(lut_f_901),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_901.INIT = 16'h8000;
LUT4 lut_inst_902 (
  .F(lut_f_902),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_902.INIT = 16'h8000;
LUT4 lut_inst_903 (
  .F(lut_f_903),
  .I0(lut_f_900),
  .I1(lut_f_901),
  .I2(lut_f_902),
  .I3(gw_vcc)
);
defparam lut_inst_903.INIT = 16'h8000;
LUT4 lut_inst_904 (
  .F(lut_f_904),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_904.INIT = 16'h8000;
LUT4 lut_inst_905 (
  .F(lut_f_905),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_905.INIT = 16'h8000;
LUT4 lut_inst_906 (
  .F(lut_f_906),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_906.INIT = 16'h8000;
LUT4 lut_inst_907 (
  .F(lut_f_907),
  .I0(lut_f_904),
  .I1(lut_f_905),
  .I2(lut_f_906),
  .I3(gw_vcc)
);
defparam lut_inst_907.INIT = 16'h8000;
LUT4 lut_inst_908 (
  .F(lut_f_908),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_908.INIT = 16'h8000;
LUT4 lut_inst_909 (
  .F(lut_f_909),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_909.INIT = 16'h8000;
LUT4 lut_inst_910 (
  .F(lut_f_910),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_910.INIT = 16'h8000;
LUT4 lut_inst_911 (
  .F(lut_f_911),
  .I0(lut_f_908),
  .I1(lut_f_909),
  .I2(lut_f_910),
  .I3(gw_vcc)
);
defparam lut_inst_911.INIT = 16'h8000;
LUT4 lut_inst_912 (
  .F(lut_f_912),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_912.INIT = 16'h8000;
LUT4 lut_inst_913 (
  .F(lut_f_913),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_913.INIT = 16'h8000;
LUT4 lut_inst_914 (
  .F(lut_f_914),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_914.INIT = 16'h8000;
LUT4 lut_inst_915 (
  .F(lut_f_915),
  .I0(lut_f_912),
  .I1(lut_f_913),
  .I2(lut_f_914),
  .I3(gw_vcc)
);
defparam lut_inst_915.INIT = 16'h8000;
LUT4 lut_inst_916 (
  .F(lut_f_916),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_916.INIT = 16'h8000;
LUT4 lut_inst_917 (
  .F(lut_f_917),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_917.INIT = 16'h8000;
LUT4 lut_inst_918 (
  .F(lut_f_918),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_918.INIT = 16'h8000;
LUT4 lut_inst_919 (
  .F(lut_f_919),
  .I0(lut_f_916),
  .I1(lut_f_917),
  .I2(lut_f_918),
  .I3(gw_vcc)
);
defparam lut_inst_919.INIT = 16'h8000;
LUT4 lut_inst_920 (
  .F(lut_f_920),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_920.INIT = 16'h8000;
LUT4 lut_inst_921 (
  .F(lut_f_921),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_921.INIT = 16'h8000;
LUT4 lut_inst_922 (
  .F(lut_f_922),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_922.INIT = 16'h8000;
LUT4 lut_inst_923 (
  .F(lut_f_923),
  .I0(lut_f_920),
  .I1(lut_f_921),
  .I2(lut_f_922),
  .I3(gw_vcc)
);
defparam lut_inst_923.INIT = 16'h8000;
LUT4 lut_inst_924 (
  .F(lut_f_924),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_924.INIT = 16'h8000;
LUT4 lut_inst_925 (
  .F(lut_f_925),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_925.INIT = 16'h8000;
LUT4 lut_inst_926 (
  .F(lut_f_926),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_926.INIT = 16'h8000;
LUT4 lut_inst_927 (
  .F(lut_f_927),
  .I0(lut_f_924),
  .I1(lut_f_925),
  .I2(lut_f_926),
  .I3(gw_vcc)
);
defparam lut_inst_927.INIT = 16'h8000;
LUT4 lut_inst_928 (
  .F(lut_f_928),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_928.INIT = 16'h8000;
LUT4 lut_inst_929 (
  .F(lut_f_929),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_929.INIT = 16'h8000;
LUT4 lut_inst_930 (
  .F(lut_f_930),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_930.INIT = 16'h8000;
LUT4 lut_inst_931 (
  .F(lut_f_931),
  .I0(lut_f_928),
  .I1(lut_f_929),
  .I2(lut_f_930),
  .I3(gw_vcc)
);
defparam lut_inst_931.INIT = 16'h8000;
LUT4 lut_inst_932 (
  .F(lut_f_932),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_932.INIT = 16'h8000;
LUT4 lut_inst_933 (
  .F(lut_f_933),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_933.INIT = 16'h8000;
LUT4 lut_inst_934 (
  .F(lut_f_934),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_934.INIT = 16'h8000;
LUT4 lut_inst_935 (
  .F(lut_f_935),
  .I0(lut_f_932),
  .I1(lut_f_933),
  .I2(lut_f_934),
  .I3(gw_vcc)
);
defparam lut_inst_935.INIT = 16'h8000;
LUT4 lut_inst_936 (
  .F(lut_f_936),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_936.INIT = 16'h8000;
LUT4 lut_inst_937 (
  .F(lut_f_937),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_937.INIT = 16'h8000;
LUT4 lut_inst_938 (
  .F(lut_f_938),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_938.INIT = 16'h8000;
LUT4 lut_inst_939 (
  .F(lut_f_939),
  .I0(lut_f_936),
  .I1(lut_f_937),
  .I2(lut_f_938),
  .I3(gw_vcc)
);
defparam lut_inst_939.INIT = 16'h8000;
LUT4 lut_inst_940 (
  .F(lut_f_940),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_940.INIT = 16'h8000;
LUT4 lut_inst_941 (
  .F(lut_f_941),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_941.INIT = 16'h8000;
LUT4 lut_inst_942 (
  .F(lut_f_942),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_942.INIT = 16'h8000;
LUT4 lut_inst_943 (
  .F(lut_f_943),
  .I0(lut_f_940),
  .I1(lut_f_941),
  .I2(lut_f_942),
  .I3(gw_vcc)
);
defparam lut_inst_943.INIT = 16'h8000;
LUT4 lut_inst_944 (
  .F(lut_f_944),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_944.INIT = 16'h8000;
LUT4 lut_inst_945 (
  .F(lut_f_945),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_945.INIT = 16'h8000;
LUT4 lut_inst_946 (
  .F(lut_f_946),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_946.INIT = 16'h8000;
LUT4 lut_inst_947 (
  .F(lut_f_947),
  .I0(lut_f_944),
  .I1(lut_f_945),
  .I2(lut_f_946),
  .I3(gw_vcc)
);
defparam lut_inst_947.INIT = 16'h8000;
LUT4 lut_inst_948 (
  .F(lut_f_948),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_948.INIT = 16'h8000;
LUT4 lut_inst_949 (
  .F(lut_f_949),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_949.INIT = 16'h8000;
LUT4 lut_inst_950 (
  .F(lut_f_950),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_950.INIT = 16'h8000;
LUT4 lut_inst_951 (
  .F(lut_f_951),
  .I0(lut_f_948),
  .I1(lut_f_949),
  .I2(lut_f_950),
  .I3(gw_vcc)
);
defparam lut_inst_951.INIT = 16'h8000;
LUT4 lut_inst_952 (
  .F(lut_f_952),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_952.INIT = 16'h8000;
LUT4 lut_inst_953 (
  .F(lut_f_953),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_953.INIT = 16'h8000;
LUT4 lut_inst_954 (
  .F(lut_f_954),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_954.INIT = 16'h8000;
LUT4 lut_inst_955 (
  .F(lut_f_955),
  .I0(lut_f_952),
  .I1(lut_f_953),
  .I2(lut_f_954),
  .I3(gw_vcc)
);
defparam lut_inst_955.INIT = 16'h8000;
LUT4 lut_inst_956 (
  .F(lut_f_956),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_956.INIT = 16'h8000;
LUT4 lut_inst_957 (
  .F(lut_f_957),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_957.INIT = 16'h8000;
LUT4 lut_inst_958 (
  .F(lut_f_958),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_958.INIT = 16'h8000;
LUT4 lut_inst_959 (
  .F(lut_f_959),
  .I0(lut_f_956),
  .I1(lut_f_957),
  .I2(lut_f_958),
  .I3(gw_vcc)
);
defparam lut_inst_959.INIT = 16'h8000;
LUT4 lut_inst_960 (
  .F(lut_f_960),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_960.INIT = 16'h8000;
LUT4 lut_inst_961 (
  .F(lut_f_961),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_961.INIT = 16'h8000;
LUT4 lut_inst_962 (
  .F(lut_f_962),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_962.INIT = 16'h8000;
LUT4 lut_inst_963 (
  .F(lut_f_963),
  .I0(lut_f_960),
  .I1(lut_f_961),
  .I2(lut_f_962),
  .I3(gw_vcc)
);
defparam lut_inst_963.INIT = 16'h8000;
LUT4 lut_inst_964 (
  .F(lut_f_964),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_964.INIT = 16'h8000;
LUT4 lut_inst_965 (
  .F(lut_f_965),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_965.INIT = 16'h8000;
LUT4 lut_inst_966 (
  .F(lut_f_966),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_966.INIT = 16'h8000;
LUT4 lut_inst_967 (
  .F(lut_f_967),
  .I0(lut_f_964),
  .I1(lut_f_965),
  .I2(lut_f_966),
  .I3(gw_vcc)
);
defparam lut_inst_967.INIT = 16'h8000;
LUT4 lut_inst_968 (
  .F(lut_f_968),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_968.INIT = 16'h8000;
LUT4 lut_inst_969 (
  .F(lut_f_969),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_969.INIT = 16'h8000;
LUT4 lut_inst_970 (
  .F(lut_f_970),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_970.INIT = 16'h8000;
LUT4 lut_inst_971 (
  .F(lut_f_971),
  .I0(lut_f_968),
  .I1(lut_f_969),
  .I2(lut_f_970),
  .I3(gw_vcc)
);
defparam lut_inst_971.INIT = 16'h8000;
LUT4 lut_inst_972 (
  .F(lut_f_972),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_972.INIT = 16'h8000;
LUT4 lut_inst_973 (
  .F(lut_f_973),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_973.INIT = 16'h8000;
LUT4 lut_inst_974 (
  .F(lut_f_974),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_974.INIT = 16'h8000;
LUT4 lut_inst_975 (
  .F(lut_f_975),
  .I0(lut_f_972),
  .I1(lut_f_973),
  .I2(lut_f_974),
  .I3(gw_vcc)
);
defparam lut_inst_975.INIT = 16'h8000;
LUT4 lut_inst_976 (
  .F(lut_f_976),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_976.INIT = 16'h8000;
LUT4 lut_inst_977 (
  .F(lut_f_977),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_977.INIT = 16'h8000;
LUT4 lut_inst_978 (
  .F(lut_f_978),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_978.INIT = 16'h8000;
LUT4 lut_inst_979 (
  .F(lut_f_979),
  .I0(lut_f_976),
  .I1(lut_f_977),
  .I2(lut_f_978),
  .I3(gw_vcc)
);
defparam lut_inst_979.INIT = 16'h8000;
LUT4 lut_inst_980 (
  .F(lut_f_980),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_980.INIT = 16'h8000;
LUT4 lut_inst_981 (
  .F(lut_f_981),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_981.INIT = 16'h8000;
LUT4 lut_inst_982 (
  .F(lut_f_982),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_982.INIT = 16'h8000;
LUT4 lut_inst_983 (
  .F(lut_f_983),
  .I0(lut_f_980),
  .I1(lut_f_981),
  .I2(lut_f_982),
  .I3(gw_vcc)
);
defparam lut_inst_983.INIT = 16'h8000;
LUT4 lut_inst_984 (
  .F(lut_f_984),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_984.INIT = 16'h8000;
LUT4 lut_inst_985 (
  .F(lut_f_985),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_985.INIT = 16'h8000;
LUT4 lut_inst_986 (
  .F(lut_f_986),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_986.INIT = 16'h8000;
LUT4 lut_inst_987 (
  .F(lut_f_987),
  .I0(lut_f_984),
  .I1(lut_f_985),
  .I2(lut_f_986),
  .I3(gw_vcc)
);
defparam lut_inst_987.INIT = 16'h8000;
LUT4 lut_inst_988 (
  .F(lut_f_988),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_988.INIT = 16'h8000;
LUT4 lut_inst_989 (
  .F(lut_f_989),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_989.INIT = 16'h8000;
LUT4 lut_inst_990 (
  .F(lut_f_990),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_990.INIT = 16'h8000;
LUT4 lut_inst_991 (
  .F(lut_f_991),
  .I0(lut_f_988),
  .I1(lut_f_989),
  .I2(lut_f_990),
  .I3(gw_vcc)
);
defparam lut_inst_991.INIT = 16'h8000;
LUT4 lut_inst_992 (
  .F(lut_f_992),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_992.INIT = 16'h8000;
LUT4 lut_inst_993 (
  .F(lut_f_993),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_993.INIT = 16'h8000;
LUT4 lut_inst_994 (
  .F(lut_f_994),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_994.INIT = 16'h8000;
LUT4 lut_inst_995 (
  .F(lut_f_995),
  .I0(lut_f_992),
  .I1(lut_f_993),
  .I2(lut_f_994),
  .I3(gw_vcc)
);
defparam lut_inst_995.INIT = 16'h8000;
LUT4 lut_inst_996 (
  .F(lut_f_996),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_996.INIT = 16'h8000;
LUT4 lut_inst_997 (
  .F(lut_f_997),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_997.INIT = 16'h8000;
LUT4 lut_inst_998 (
  .F(lut_f_998),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_998.INIT = 16'h8000;
LUT4 lut_inst_999 (
  .F(lut_f_999),
  .I0(lut_f_996),
  .I1(lut_f_997),
  .I2(lut_f_998),
  .I3(gw_vcc)
);
defparam lut_inst_999.INIT = 16'h8000;
LUT4 lut_inst_1000 (
  .F(lut_f_1000),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1000.INIT = 16'h8000;
LUT4 lut_inst_1001 (
  .F(lut_f_1001),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1001.INIT = 16'h8000;
LUT4 lut_inst_1002 (
  .F(lut_f_1002),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1002.INIT = 16'h8000;
LUT4 lut_inst_1003 (
  .F(lut_f_1003),
  .I0(lut_f_1000),
  .I1(lut_f_1001),
  .I2(lut_f_1002),
  .I3(gw_vcc)
);
defparam lut_inst_1003.INIT = 16'h8000;
LUT4 lut_inst_1004 (
  .F(lut_f_1004),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1004.INIT = 16'h8000;
LUT4 lut_inst_1005 (
  .F(lut_f_1005),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1005.INIT = 16'h8000;
LUT4 lut_inst_1006 (
  .F(lut_f_1006),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1006.INIT = 16'h8000;
LUT4 lut_inst_1007 (
  .F(lut_f_1007),
  .I0(lut_f_1004),
  .I1(lut_f_1005),
  .I2(lut_f_1006),
  .I3(gw_vcc)
);
defparam lut_inst_1007.INIT = 16'h8000;
LUT4 lut_inst_1008 (
  .F(lut_f_1008),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1008.INIT = 16'h8000;
LUT4 lut_inst_1009 (
  .F(lut_f_1009),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1009.INIT = 16'h8000;
LUT4 lut_inst_1010 (
  .F(lut_f_1010),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1010.INIT = 16'h8000;
LUT4 lut_inst_1011 (
  .F(lut_f_1011),
  .I0(lut_f_1008),
  .I1(lut_f_1009),
  .I2(lut_f_1010),
  .I3(gw_vcc)
);
defparam lut_inst_1011.INIT = 16'h8000;
LUT4 lut_inst_1012 (
  .F(lut_f_1012),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1012.INIT = 16'h8000;
LUT4 lut_inst_1013 (
  .F(lut_f_1013),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1013.INIT = 16'h8000;
LUT4 lut_inst_1014 (
  .F(lut_f_1014),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1014.INIT = 16'h8000;
LUT4 lut_inst_1015 (
  .F(lut_f_1015),
  .I0(lut_f_1012),
  .I1(lut_f_1013),
  .I2(lut_f_1014),
  .I3(gw_vcc)
);
defparam lut_inst_1015.INIT = 16'h8000;
LUT4 lut_inst_1016 (
  .F(lut_f_1016),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1016.INIT = 16'h8000;
LUT4 lut_inst_1017 (
  .F(lut_f_1017),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1017.INIT = 16'h8000;
LUT4 lut_inst_1018 (
  .F(lut_f_1018),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1018.INIT = 16'h8000;
LUT4 lut_inst_1019 (
  .F(lut_f_1019),
  .I0(lut_f_1016),
  .I1(lut_f_1017),
  .I2(lut_f_1018),
  .I3(gw_vcc)
);
defparam lut_inst_1019.INIT = 16'h8000;
LUT4 lut_inst_1020 (
  .F(lut_f_1020),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1020.INIT = 16'h8000;
LUT4 lut_inst_1021 (
  .F(lut_f_1021),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1021.INIT = 16'h8000;
LUT4 lut_inst_1022 (
  .F(lut_f_1022),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1022.INIT = 16'h8000;
LUT4 lut_inst_1023 (
  .F(lut_f_1023),
  .I0(lut_f_1020),
  .I1(lut_f_1021),
  .I2(lut_f_1022),
  .I3(gw_vcc)
);
defparam lut_inst_1023.INIT = 16'h8000;
LUT4 lut_inst_1024 (
  .F(lut_f_1024),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1024.INIT = 16'h8000;
LUT4 lut_inst_1025 (
  .F(lut_f_1025),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1025.INIT = 16'h8000;
LUT4 lut_inst_1026 (
  .F(lut_f_1026),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1026.INIT = 16'h8000;
LUT4 lut_inst_1027 (
  .F(lut_f_1027),
  .I0(lut_f_1024),
  .I1(lut_f_1025),
  .I2(lut_f_1026),
  .I3(gw_vcc)
);
defparam lut_inst_1027.INIT = 16'h8000;
LUT4 lut_inst_1028 (
  .F(lut_f_1028),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1028.INIT = 16'h8000;
LUT4 lut_inst_1029 (
  .F(lut_f_1029),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1029.INIT = 16'h8000;
LUT4 lut_inst_1030 (
  .F(lut_f_1030),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1030.INIT = 16'h8000;
LUT4 lut_inst_1031 (
  .F(lut_f_1031),
  .I0(lut_f_1028),
  .I1(lut_f_1029),
  .I2(lut_f_1030),
  .I3(gw_vcc)
);
defparam lut_inst_1031.INIT = 16'h8000;
LUT4 lut_inst_1032 (
  .F(lut_f_1032),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1032.INIT = 16'h8000;
LUT4 lut_inst_1033 (
  .F(lut_f_1033),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1033.INIT = 16'h8000;
LUT4 lut_inst_1034 (
  .F(lut_f_1034),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1034.INIT = 16'h8000;
LUT4 lut_inst_1035 (
  .F(lut_f_1035),
  .I0(lut_f_1032),
  .I1(lut_f_1033),
  .I2(lut_f_1034),
  .I3(gw_vcc)
);
defparam lut_inst_1035.INIT = 16'h8000;
LUT4 lut_inst_1036 (
  .F(lut_f_1036),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1036.INIT = 16'h8000;
LUT4 lut_inst_1037 (
  .F(lut_f_1037),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1037.INIT = 16'h8000;
LUT4 lut_inst_1038 (
  .F(lut_f_1038),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1038.INIT = 16'h8000;
LUT4 lut_inst_1039 (
  .F(lut_f_1039),
  .I0(lut_f_1036),
  .I1(lut_f_1037),
  .I2(lut_f_1038),
  .I3(gw_vcc)
);
defparam lut_inst_1039.INIT = 16'h8000;
LUT4 lut_inst_1040 (
  .F(lut_f_1040),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1040.INIT = 16'h8000;
LUT4 lut_inst_1041 (
  .F(lut_f_1041),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1041.INIT = 16'h8000;
LUT4 lut_inst_1042 (
  .F(lut_f_1042),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1042.INIT = 16'h8000;
LUT4 lut_inst_1043 (
  .F(lut_f_1043),
  .I0(lut_f_1040),
  .I1(lut_f_1041),
  .I2(lut_f_1042),
  .I3(gw_vcc)
);
defparam lut_inst_1043.INIT = 16'h8000;
LUT4 lut_inst_1044 (
  .F(lut_f_1044),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1044.INIT = 16'h8000;
LUT4 lut_inst_1045 (
  .F(lut_f_1045),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1045.INIT = 16'h8000;
LUT4 lut_inst_1046 (
  .F(lut_f_1046),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1046.INIT = 16'h8000;
LUT4 lut_inst_1047 (
  .F(lut_f_1047),
  .I0(lut_f_1044),
  .I1(lut_f_1045),
  .I2(lut_f_1046),
  .I3(gw_vcc)
);
defparam lut_inst_1047.INIT = 16'h8000;
LUT4 lut_inst_1048 (
  .F(lut_f_1048),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1048.INIT = 16'h8000;
LUT4 lut_inst_1049 (
  .F(lut_f_1049),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1049.INIT = 16'h8000;
LUT4 lut_inst_1050 (
  .F(lut_f_1050),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1050.INIT = 16'h8000;
LUT4 lut_inst_1051 (
  .F(lut_f_1051),
  .I0(lut_f_1048),
  .I1(lut_f_1049),
  .I2(lut_f_1050),
  .I3(gw_vcc)
);
defparam lut_inst_1051.INIT = 16'h8000;
LUT4 lut_inst_1052 (
  .F(lut_f_1052),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1052.INIT = 16'h8000;
LUT4 lut_inst_1053 (
  .F(lut_f_1053),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1053.INIT = 16'h8000;
LUT4 lut_inst_1054 (
  .F(lut_f_1054),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1054.INIT = 16'h8000;
LUT4 lut_inst_1055 (
  .F(lut_f_1055),
  .I0(lut_f_1052),
  .I1(lut_f_1053),
  .I2(lut_f_1054),
  .I3(gw_vcc)
);
defparam lut_inst_1055.INIT = 16'h8000;
LUT4 lut_inst_1056 (
  .F(lut_f_1056),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1056.INIT = 16'h8000;
LUT4 lut_inst_1057 (
  .F(lut_f_1057),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1057.INIT = 16'h8000;
LUT4 lut_inst_1058 (
  .F(lut_f_1058),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1058.INIT = 16'h8000;
LUT4 lut_inst_1059 (
  .F(lut_f_1059),
  .I0(lut_f_1056),
  .I1(lut_f_1057),
  .I2(lut_f_1058),
  .I3(gw_vcc)
);
defparam lut_inst_1059.INIT = 16'h8000;
LUT4 lut_inst_1060 (
  .F(lut_f_1060),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1060.INIT = 16'h8000;
LUT4 lut_inst_1061 (
  .F(lut_f_1061),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1061.INIT = 16'h8000;
LUT4 lut_inst_1062 (
  .F(lut_f_1062),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1062.INIT = 16'h8000;
LUT4 lut_inst_1063 (
  .F(lut_f_1063),
  .I0(lut_f_1060),
  .I1(lut_f_1061),
  .I2(lut_f_1062),
  .I3(gw_vcc)
);
defparam lut_inst_1063.INIT = 16'h8000;
LUT4 lut_inst_1064 (
  .F(lut_f_1064),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1064.INIT = 16'h8000;
LUT4 lut_inst_1065 (
  .F(lut_f_1065),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1065.INIT = 16'h8000;
LUT4 lut_inst_1066 (
  .F(lut_f_1066),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1066.INIT = 16'h8000;
LUT4 lut_inst_1067 (
  .F(lut_f_1067),
  .I0(lut_f_1064),
  .I1(lut_f_1065),
  .I2(lut_f_1066),
  .I3(gw_vcc)
);
defparam lut_inst_1067.INIT = 16'h8000;
LUT4 lut_inst_1068 (
  .F(lut_f_1068),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1068.INIT = 16'h8000;
LUT4 lut_inst_1069 (
  .F(lut_f_1069),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1069.INIT = 16'h8000;
LUT4 lut_inst_1070 (
  .F(lut_f_1070),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1070.INIT = 16'h8000;
LUT4 lut_inst_1071 (
  .F(lut_f_1071),
  .I0(lut_f_1068),
  .I1(lut_f_1069),
  .I2(lut_f_1070),
  .I3(gw_vcc)
);
defparam lut_inst_1071.INIT = 16'h8000;
LUT4 lut_inst_1072 (
  .F(lut_f_1072),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1072.INIT = 16'h8000;
LUT4 lut_inst_1073 (
  .F(lut_f_1073),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1073.INIT = 16'h8000;
LUT4 lut_inst_1074 (
  .F(lut_f_1074),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1074.INIT = 16'h8000;
LUT4 lut_inst_1075 (
  .F(lut_f_1075),
  .I0(lut_f_1072),
  .I1(lut_f_1073),
  .I2(lut_f_1074),
  .I3(gw_vcc)
);
defparam lut_inst_1075.INIT = 16'h8000;
LUT4 lut_inst_1076 (
  .F(lut_f_1076),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1076.INIT = 16'h8000;
LUT4 lut_inst_1077 (
  .F(lut_f_1077),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1077.INIT = 16'h8000;
LUT4 lut_inst_1078 (
  .F(lut_f_1078),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1078.INIT = 16'h8000;
LUT4 lut_inst_1079 (
  .F(lut_f_1079),
  .I0(lut_f_1076),
  .I1(lut_f_1077),
  .I2(lut_f_1078),
  .I3(gw_vcc)
);
defparam lut_inst_1079.INIT = 16'h8000;
LUT4 lut_inst_1080 (
  .F(lut_f_1080),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1080.INIT = 16'h8000;
LUT4 lut_inst_1081 (
  .F(lut_f_1081),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1081.INIT = 16'h8000;
LUT4 lut_inst_1082 (
  .F(lut_f_1082),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1082.INIT = 16'h8000;
LUT4 lut_inst_1083 (
  .F(lut_f_1083),
  .I0(lut_f_1080),
  .I1(lut_f_1081),
  .I2(lut_f_1082),
  .I3(gw_vcc)
);
defparam lut_inst_1083.INIT = 16'h8000;
LUT4 lut_inst_1084 (
  .F(lut_f_1084),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1084.INIT = 16'h8000;
LUT4 lut_inst_1085 (
  .F(lut_f_1085),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1085.INIT = 16'h8000;
LUT4 lut_inst_1086 (
  .F(lut_f_1086),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1086.INIT = 16'h8000;
LUT4 lut_inst_1087 (
  .F(lut_f_1087),
  .I0(lut_f_1084),
  .I1(lut_f_1085),
  .I2(lut_f_1086),
  .I3(gw_vcc)
);
defparam lut_inst_1087.INIT = 16'h8000;
LUT4 lut_inst_1088 (
  .F(lut_f_1088),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1088.INIT = 16'h8000;
LUT4 lut_inst_1089 (
  .F(lut_f_1089),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1089.INIT = 16'h8000;
LUT4 lut_inst_1090 (
  .F(lut_f_1090),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1090.INIT = 16'h8000;
LUT4 lut_inst_1091 (
  .F(lut_f_1091),
  .I0(lut_f_1088),
  .I1(lut_f_1089),
  .I2(lut_f_1090),
  .I3(gw_vcc)
);
defparam lut_inst_1091.INIT = 16'h8000;
LUT4 lut_inst_1092 (
  .F(lut_f_1092),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1092.INIT = 16'h8000;
LUT4 lut_inst_1093 (
  .F(lut_f_1093),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1093.INIT = 16'h8000;
LUT4 lut_inst_1094 (
  .F(lut_f_1094),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1094.INIT = 16'h8000;
LUT4 lut_inst_1095 (
  .F(lut_f_1095),
  .I0(lut_f_1092),
  .I1(lut_f_1093),
  .I2(lut_f_1094),
  .I3(gw_vcc)
);
defparam lut_inst_1095.INIT = 16'h8000;
LUT4 lut_inst_1096 (
  .F(lut_f_1096),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1096.INIT = 16'h8000;
LUT4 lut_inst_1097 (
  .F(lut_f_1097),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1097.INIT = 16'h8000;
LUT4 lut_inst_1098 (
  .F(lut_f_1098),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1098.INIT = 16'h8000;
LUT4 lut_inst_1099 (
  .F(lut_f_1099),
  .I0(lut_f_1096),
  .I1(lut_f_1097),
  .I2(lut_f_1098),
  .I3(gw_vcc)
);
defparam lut_inst_1099.INIT = 16'h8000;
LUT4 lut_inst_1100 (
  .F(lut_f_1100),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1100.INIT = 16'h8000;
LUT4 lut_inst_1101 (
  .F(lut_f_1101),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1101.INIT = 16'h8000;
LUT4 lut_inst_1102 (
  .F(lut_f_1102),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1102.INIT = 16'h8000;
LUT4 lut_inst_1103 (
  .F(lut_f_1103),
  .I0(lut_f_1100),
  .I1(lut_f_1101),
  .I2(lut_f_1102),
  .I3(gw_vcc)
);
defparam lut_inst_1103.INIT = 16'h8000;
LUT4 lut_inst_1104 (
  .F(lut_f_1104),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1104.INIT = 16'h8000;
LUT4 lut_inst_1105 (
  .F(lut_f_1105),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1105.INIT = 16'h8000;
LUT4 lut_inst_1106 (
  .F(lut_f_1106),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1106.INIT = 16'h8000;
LUT4 lut_inst_1107 (
  .F(lut_f_1107),
  .I0(lut_f_1104),
  .I1(lut_f_1105),
  .I2(lut_f_1106),
  .I3(gw_vcc)
);
defparam lut_inst_1107.INIT = 16'h8000;
LUT4 lut_inst_1108 (
  .F(lut_f_1108),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1108.INIT = 16'h8000;
LUT4 lut_inst_1109 (
  .F(lut_f_1109),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1109.INIT = 16'h8000;
LUT4 lut_inst_1110 (
  .F(lut_f_1110),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1110.INIT = 16'h8000;
LUT4 lut_inst_1111 (
  .F(lut_f_1111),
  .I0(lut_f_1108),
  .I1(lut_f_1109),
  .I2(lut_f_1110),
  .I3(gw_vcc)
);
defparam lut_inst_1111.INIT = 16'h8000;
LUT4 lut_inst_1112 (
  .F(lut_f_1112),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1112.INIT = 16'h8000;
LUT4 lut_inst_1113 (
  .F(lut_f_1113),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1113.INIT = 16'h8000;
LUT4 lut_inst_1114 (
  .F(lut_f_1114),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1114.INIT = 16'h8000;
LUT4 lut_inst_1115 (
  .F(lut_f_1115),
  .I0(lut_f_1112),
  .I1(lut_f_1113),
  .I2(lut_f_1114),
  .I3(gw_vcc)
);
defparam lut_inst_1115.INIT = 16'h8000;
LUT4 lut_inst_1116 (
  .F(lut_f_1116),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1116.INIT = 16'h8000;
LUT4 lut_inst_1117 (
  .F(lut_f_1117),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1117.INIT = 16'h8000;
LUT4 lut_inst_1118 (
  .F(lut_f_1118),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1118.INIT = 16'h8000;
LUT4 lut_inst_1119 (
  .F(lut_f_1119),
  .I0(lut_f_1116),
  .I1(lut_f_1117),
  .I2(lut_f_1118),
  .I3(gw_vcc)
);
defparam lut_inst_1119.INIT = 16'h8000;
LUT4 lut_inst_1120 (
  .F(lut_f_1120),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1120.INIT = 16'h8000;
LUT4 lut_inst_1121 (
  .F(lut_f_1121),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1121.INIT = 16'h8000;
LUT4 lut_inst_1122 (
  .F(lut_f_1122),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1122.INIT = 16'h8000;
LUT4 lut_inst_1123 (
  .F(lut_f_1123),
  .I0(lut_f_1120),
  .I1(lut_f_1121),
  .I2(lut_f_1122),
  .I3(gw_vcc)
);
defparam lut_inst_1123.INIT = 16'h8000;
LUT4 lut_inst_1124 (
  .F(lut_f_1124),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1124.INIT = 16'h8000;
LUT4 lut_inst_1125 (
  .F(lut_f_1125),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1125.INIT = 16'h8000;
LUT4 lut_inst_1126 (
  .F(lut_f_1126),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1126.INIT = 16'h8000;
LUT4 lut_inst_1127 (
  .F(lut_f_1127),
  .I0(lut_f_1124),
  .I1(lut_f_1125),
  .I2(lut_f_1126),
  .I3(gw_vcc)
);
defparam lut_inst_1127.INIT = 16'h8000;
LUT4 lut_inst_1128 (
  .F(lut_f_1128),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1128.INIT = 16'h8000;
LUT4 lut_inst_1129 (
  .F(lut_f_1129),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1129.INIT = 16'h8000;
LUT4 lut_inst_1130 (
  .F(lut_f_1130),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1130.INIT = 16'h8000;
LUT4 lut_inst_1131 (
  .F(lut_f_1131),
  .I0(lut_f_1128),
  .I1(lut_f_1129),
  .I2(lut_f_1130),
  .I3(gw_vcc)
);
defparam lut_inst_1131.INIT = 16'h8000;
LUT4 lut_inst_1132 (
  .F(lut_f_1132),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1132.INIT = 16'h8000;
LUT4 lut_inst_1133 (
  .F(lut_f_1133),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1133.INIT = 16'h8000;
LUT4 lut_inst_1134 (
  .F(lut_f_1134),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1134.INIT = 16'h8000;
LUT4 lut_inst_1135 (
  .F(lut_f_1135),
  .I0(lut_f_1132),
  .I1(lut_f_1133),
  .I2(lut_f_1134),
  .I3(gw_vcc)
);
defparam lut_inst_1135.INIT = 16'h8000;
LUT4 lut_inst_1136 (
  .F(lut_f_1136),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1136.INIT = 16'h8000;
LUT4 lut_inst_1137 (
  .F(lut_f_1137),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1137.INIT = 16'h8000;
LUT4 lut_inst_1138 (
  .F(lut_f_1138),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1138.INIT = 16'h8000;
LUT4 lut_inst_1139 (
  .F(lut_f_1139),
  .I0(lut_f_1136),
  .I1(lut_f_1137),
  .I2(lut_f_1138),
  .I3(gw_vcc)
);
defparam lut_inst_1139.INIT = 16'h8000;
LUT4 lut_inst_1140 (
  .F(lut_f_1140),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1140.INIT = 16'h8000;
LUT4 lut_inst_1141 (
  .F(lut_f_1141),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1141.INIT = 16'h8000;
LUT4 lut_inst_1142 (
  .F(lut_f_1142),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1142.INIT = 16'h8000;
LUT4 lut_inst_1143 (
  .F(lut_f_1143),
  .I0(lut_f_1140),
  .I1(lut_f_1141),
  .I2(lut_f_1142),
  .I3(gw_vcc)
);
defparam lut_inst_1143.INIT = 16'h8000;
LUT4 lut_inst_1144 (
  .F(lut_f_1144),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1144.INIT = 16'h8000;
LUT4 lut_inst_1145 (
  .F(lut_f_1145),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1145.INIT = 16'h8000;
LUT4 lut_inst_1146 (
  .F(lut_f_1146),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1146.INIT = 16'h8000;
LUT4 lut_inst_1147 (
  .F(lut_f_1147),
  .I0(lut_f_1144),
  .I1(lut_f_1145),
  .I2(lut_f_1146),
  .I3(gw_vcc)
);
defparam lut_inst_1147.INIT = 16'h8000;
LUT4 lut_inst_1148 (
  .F(lut_f_1148),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1148.INIT = 16'h8000;
LUT4 lut_inst_1149 (
  .F(lut_f_1149),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1149.INIT = 16'h8000;
LUT4 lut_inst_1150 (
  .F(lut_f_1150),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1150.INIT = 16'h8000;
LUT4 lut_inst_1151 (
  .F(lut_f_1151),
  .I0(lut_f_1148),
  .I1(lut_f_1149),
  .I2(lut_f_1150),
  .I3(gw_vcc)
);
defparam lut_inst_1151.INIT = 16'h8000;
LUT4 lut_inst_1152 (
  .F(lut_f_1152),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1152.INIT = 16'h8000;
LUT4 lut_inst_1153 (
  .F(lut_f_1153),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1153.INIT = 16'h8000;
LUT4 lut_inst_1154 (
  .F(lut_f_1154),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1154.INIT = 16'h8000;
LUT4 lut_inst_1155 (
  .F(lut_f_1155),
  .I0(lut_f_1152),
  .I1(lut_f_1153),
  .I2(lut_f_1154),
  .I3(gw_vcc)
);
defparam lut_inst_1155.INIT = 16'h8000;
LUT4 lut_inst_1156 (
  .F(lut_f_1156),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1156.INIT = 16'h8000;
LUT4 lut_inst_1157 (
  .F(lut_f_1157),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1157.INIT = 16'h8000;
LUT4 lut_inst_1158 (
  .F(lut_f_1158),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1158.INIT = 16'h8000;
LUT4 lut_inst_1159 (
  .F(lut_f_1159),
  .I0(lut_f_1156),
  .I1(lut_f_1157),
  .I2(lut_f_1158),
  .I3(gw_vcc)
);
defparam lut_inst_1159.INIT = 16'h8000;
LUT4 lut_inst_1160 (
  .F(lut_f_1160),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1160.INIT = 16'h8000;
LUT4 lut_inst_1161 (
  .F(lut_f_1161),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1161.INIT = 16'h8000;
LUT4 lut_inst_1162 (
  .F(lut_f_1162),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1162.INIT = 16'h8000;
LUT4 lut_inst_1163 (
  .F(lut_f_1163),
  .I0(lut_f_1160),
  .I1(lut_f_1161),
  .I2(lut_f_1162),
  .I3(gw_vcc)
);
defparam lut_inst_1163.INIT = 16'h8000;
LUT4 lut_inst_1164 (
  .F(lut_f_1164),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1164.INIT = 16'h8000;
LUT4 lut_inst_1165 (
  .F(lut_f_1165),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1165.INIT = 16'h8000;
LUT4 lut_inst_1166 (
  .F(lut_f_1166),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1166.INIT = 16'h8000;
LUT4 lut_inst_1167 (
  .F(lut_f_1167),
  .I0(lut_f_1164),
  .I1(lut_f_1165),
  .I2(lut_f_1166),
  .I3(gw_vcc)
);
defparam lut_inst_1167.INIT = 16'h8000;
LUT4 lut_inst_1168 (
  .F(lut_f_1168),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1168.INIT = 16'h8000;
LUT4 lut_inst_1169 (
  .F(lut_f_1169),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1169.INIT = 16'h8000;
LUT4 lut_inst_1170 (
  .F(lut_f_1170),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1170.INIT = 16'h8000;
LUT4 lut_inst_1171 (
  .F(lut_f_1171),
  .I0(lut_f_1168),
  .I1(lut_f_1169),
  .I2(lut_f_1170),
  .I3(gw_vcc)
);
defparam lut_inst_1171.INIT = 16'h8000;
LUT4 lut_inst_1172 (
  .F(lut_f_1172),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1172.INIT = 16'h8000;
LUT4 lut_inst_1173 (
  .F(lut_f_1173),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1173.INIT = 16'h8000;
LUT4 lut_inst_1174 (
  .F(lut_f_1174),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1174.INIT = 16'h8000;
LUT4 lut_inst_1175 (
  .F(lut_f_1175),
  .I0(lut_f_1172),
  .I1(lut_f_1173),
  .I2(lut_f_1174),
  .I3(gw_vcc)
);
defparam lut_inst_1175.INIT = 16'h8000;
LUT4 lut_inst_1176 (
  .F(lut_f_1176),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1176.INIT = 16'h8000;
LUT4 lut_inst_1177 (
  .F(lut_f_1177),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1177.INIT = 16'h8000;
LUT4 lut_inst_1178 (
  .F(lut_f_1178),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1178.INIT = 16'h8000;
LUT4 lut_inst_1179 (
  .F(lut_f_1179),
  .I0(lut_f_1176),
  .I1(lut_f_1177),
  .I2(lut_f_1178),
  .I3(gw_vcc)
);
defparam lut_inst_1179.INIT = 16'h8000;
LUT4 lut_inst_1180 (
  .F(lut_f_1180),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1180.INIT = 16'h8000;
LUT4 lut_inst_1181 (
  .F(lut_f_1181),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1181.INIT = 16'h8000;
LUT4 lut_inst_1182 (
  .F(lut_f_1182),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1182.INIT = 16'h8000;
LUT4 lut_inst_1183 (
  .F(lut_f_1183),
  .I0(lut_f_1180),
  .I1(lut_f_1181),
  .I2(lut_f_1182),
  .I3(gw_vcc)
);
defparam lut_inst_1183.INIT = 16'h8000;
LUT4 lut_inst_1184 (
  .F(lut_f_1184),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1184.INIT = 16'h8000;
LUT4 lut_inst_1185 (
  .F(lut_f_1185),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1185.INIT = 16'h8000;
LUT4 lut_inst_1186 (
  .F(lut_f_1186),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1186.INIT = 16'h8000;
LUT4 lut_inst_1187 (
  .F(lut_f_1187),
  .I0(lut_f_1184),
  .I1(lut_f_1185),
  .I2(lut_f_1186),
  .I3(gw_vcc)
);
defparam lut_inst_1187.INIT = 16'h8000;
LUT4 lut_inst_1188 (
  .F(lut_f_1188),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1188.INIT = 16'h8000;
LUT4 lut_inst_1189 (
  .F(lut_f_1189),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1189.INIT = 16'h8000;
LUT4 lut_inst_1190 (
  .F(lut_f_1190),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1190.INIT = 16'h8000;
LUT4 lut_inst_1191 (
  .F(lut_f_1191),
  .I0(lut_f_1188),
  .I1(lut_f_1189),
  .I2(lut_f_1190),
  .I3(gw_vcc)
);
defparam lut_inst_1191.INIT = 16'h8000;
LUT4 lut_inst_1192 (
  .F(lut_f_1192),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1192.INIT = 16'h8000;
LUT4 lut_inst_1193 (
  .F(lut_f_1193),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1193.INIT = 16'h8000;
LUT4 lut_inst_1194 (
  .F(lut_f_1194),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1194.INIT = 16'h8000;
LUT4 lut_inst_1195 (
  .F(lut_f_1195),
  .I0(lut_f_1192),
  .I1(lut_f_1193),
  .I2(lut_f_1194),
  .I3(gw_vcc)
);
defparam lut_inst_1195.INIT = 16'h8000;
LUT4 lut_inst_1196 (
  .F(lut_f_1196),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1196.INIT = 16'h8000;
LUT4 lut_inst_1197 (
  .F(lut_f_1197),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1197.INIT = 16'h8000;
LUT4 lut_inst_1198 (
  .F(lut_f_1198),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1198.INIT = 16'h8000;
LUT4 lut_inst_1199 (
  .F(lut_f_1199),
  .I0(lut_f_1196),
  .I1(lut_f_1197),
  .I2(lut_f_1198),
  .I3(gw_vcc)
);
defparam lut_inst_1199.INIT = 16'h8000;
LUT4 lut_inst_1200 (
  .F(lut_f_1200),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1200.INIT = 16'h8000;
LUT4 lut_inst_1201 (
  .F(lut_f_1201),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1201.INIT = 16'h8000;
LUT4 lut_inst_1202 (
  .F(lut_f_1202),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1202.INIT = 16'h8000;
LUT4 lut_inst_1203 (
  .F(lut_f_1203),
  .I0(lut_f_1200),
  .I1(lut_f_1201),
  .I2(lut_f_1202),
  .I3(gw_vcc)
);
defparam lut_inst_1203.INIT = 16'h8000;
LUT4 lut_inst_1204 (
  .F(lut_f_1204),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1204.INIT = 16'h8000;
LUT4 lut_inst_1205 (
  .F(lut_f_1205),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1205.INIT = 16'h8000;
LUT4 lut_inst_1206 (
  .F(lut_f_1206),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1206.INIT = 16'h8000;
LUT4 lut_inst_1207 (
  .F(lut_f_1207),
  .I0(lut_f_1204),
  .I1(lut_f_1205),
  .I2(lut_f_1206),
  .I3(gw_vcc)
);
defparam lut_inst_1207.INIT = 16'h8000;
LUT4 lut_inst_1208 (
  .F(lut_f_1208),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1208.INIT = 16'h8000;
LUT4 lut_inst_1209 (
  .F(lut_f_1209),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1209.INIT = 16'h8000;
LUT4 lut_inst_1210 (
  .F(lut_f_1210),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1210.INIT = 16'h8000;
LUT4 lut_inst_1211 (
  .F(lut_f_1211),
  .I0(lut_f_1208),
  .I1(lut_f_1209),
  .I2(lut_f_1210),
  .I3(gw_vcc)
);
defparam lut_inst_1211.INIT = 16'h8000;
LUT4 lut_inst_1212 (
  .F(lut_f_1212),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1212.INIT = 16'h8000;
LUT4 lut_inst_1213 (
  .F(lut_f_1213),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1213.INIT = 16'h8000;
LUT4 lut_inst_1214 (
  .F(lut_f_1214),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1214.INIT = 16'h8000;
LUT4 lut_inst_1215 (
  .F(lut_f_1215),
  .I0(lut_f_1212),
  .I1(lut_f_1213),
  .I2(lut_f_1214),
  .I3(gw_vcc)
);
defparam lut_inst_1215.INIT = 16'h8000;
LUT4 lut_inst_1216 (
  .F(lut_f_1216),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1216.INIT = 16'h8000;
LUT4 lut_inst_1217 (
  .F(lut_f_1217),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1217.INIT = 16'h8000;
LUT4 lut_inst_1218 (
  .F(lut_f_1218),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1218.INIT = 16'h8000;
LUT4 lut_inst_1219 (
  .F(lut_f_1219),
  .I0(lut_f_1216),
  .I1(lut_f_1217),
  .I2(lut_f_1218),
  .I3(gw_vcc)
);
defparam lut_inst_1219.INIT = 16'h8000;
LUT4 lut_inst_1220 (
  .F(lut_f_1220),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1220.INIT = 16'h8000;
LUT4 lut_inst_1221 (
  .F(lut_f_1221),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1221.INIT = 16'h8000;
LUT4 lut_inst_1222 (
  .F(lut_f_1222),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1222.INIT = 16'h8000;
LUT4 lut_inst_1223 (
  .F(lut_f_1223),
  .I0(lut_f_1220),
  .I1(lut_f_1221),
  .I2(lut_f_1222),
  .I3(gw_vcc)
);
defparam lut_inst_1223.INIT = 16'h8000;
LUT4 lut_inst_1224 (
  .F(lut_f_1224),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1224.INIT = 16'h8000;
LUT4 lut_inst_1225 (
  .F(lut_f_1225),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1225.INIT = 16'h8000;
LUT4 lut_inst_1226 (
  .F(lut_f_1226),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1226.INIT = 16'h8000;
LUT4 lut_inst_1227 (
  .F(lut_f_1227),
  .I0(lut_f_1224),
  .I1(lut_f_1225),
  .I2(lut_f_1226),
  .I3(gw_vcc)
);
defparam lut_inst_1227.INIT = 16'h8000;
LUT4 lut_inst_1228 (
  .F(lut_f_1228),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1228.INIT = 16'h8000;
LUT4 lut_inst_1229 (
  .F(lut_f_1229),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1229.INIT = 16'h8000;
LUT4 lut_inst_1230 (
  .F(lut_f_1230),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1230.INIT = 16'h8000;
LUT4 lut_inst_1231 (
  .F(lut_f_1231),
  .I0(lut_f_1228),
  .I1(lut_f_1229),
  .I2(lut_f_1230),
  .I3(gw_vcc)
);
defparam lut_inst_1231.INIT = 16'h8000;
LUT4 lut_inst_1232 (
  .F(lut_f_1232),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1232.INIT = 16'h8000;
LUT4 lut_inst_1233 (
  .F(lut_f_1233),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1233.INIT = 16'h8000;
LUT4 lut_inst_1234 (
  .F(lut_f_1234),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1234.INIT = 16'h8000;
LUT4 lut_inst_1235 (
  .F(lut_f_1235),
  .I0(lut_f_1232),
  .I1(lut_f_1233),
  .I2(lut_f_1234),
  .I3(gw_vcc)
);
defparam lut_inst_1235.INIT = 16'h8000;
LUT4 lut_inst_1236 (
  .F(lut_f_1236),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1236.INIT = 16'h8000;
LUT4 lut_inst_1237 (
  .F(lut_f_1237),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1237.INIT = 16'h8000;
LUT4 lut_inst_1238 (
  .F(lut_f_1238),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1238.INIT = 16'h8000;
LUT4 lut_inst_1239 (
  .F(lut_f_1239),
  .I0(lut_f_1236),
  .I1(lut_f_1237),
  .I2(lut_f_1238),
  .I3(gw_vcc)
);
defparam lut_inst_1239.INIT = 16'h8000;
LUT4 lut_inst_1240 (
  .F(lut_f_1240),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1240.INIT = 16'h8000;
LUT4 lut_inst_1241 (
  .F(lut_f_1241),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1241.INIT = 16'h8000;
LUT4 lut_inst_1242 (
  .F(lut_f_1242),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1242.INIT = 16'h8000;
LUT4 lut_inst_1243 (
  .F(lut_f_1243),
  .I0(lut_f_1240),
  .I1(lut_f_1241),
  .I2(lut_f_1242),
  .I3(gw_vcc)
);
defparam lut_inst_1243.INIT = 16'h8000;
LUT4 lut_inst_1244 (
  .F(lut_f_1244),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1244.INIT = 16'h8000;
LUT4 lut_inst_1245 (
  .F(lut_f_1245),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1245.INIT = 16'h8000;
LUT4 lut_inst_1246 (
  .F(lut_f_1246),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1246.INIT = 16'h8000;
LUT4 lut_inst_1247 (
  .F(lut_f_1247),
  .I0(lut_f_1244),
  .I1(lut_f_1245),
  .I2(lut_f_1246),
  .I3(gw_vcc)
);
defparam lut_inst_1247.INIT = 16'h8000;
LUT4 lut_inst_1248 (
  .F(lut_f_1248),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1248.INIT = 16'h8000;
LUT4 lut_inst_1249 (
  .F(lut_f_1249),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1249.INIT = 16'h8000;
LUT4 lut_inst_1250 (
  .F(lut_f_1250),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1250.INIT = 16'h8000;
LUT4 lut_inst_1251 (
  .F(lut_f_1251),
  .I0(lut_f_1248),
  .I1(lut_f_1249),
  .I2(lut_f_1250),
  .I3(gw_vcc)
);
defparam lut_inst_1251.INIT = 16'h8000;
LUT4 lut_inst_1252 (
  .F(lut_f_1252),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1252.INIT = 16'h8000;
LUT4 lut_inst_1253 (
  .F(lut_f_1253),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1253.INIT = 16'h8000;
LUT4 lut_inst_1254 (
  .F(lut_f_1254),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1254.INIT = 16'h8000;
LUT4 lut_inst_1255 (
  .F(lut_f_1255),
  .I0(lut_f_1252),
  .I1(lut_f_1253),
  .I2(lut_f_1254),
  .I3(gw_vcc)
);
defparam lut_inst_1255.INIT = 16'h8000;
LUT4 lut_inst_1256 (
  .F(lut_f_1256),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1256.INIT = 16'h8000;
LUT4 lut_inst_1257 (
  .F(lut_f_1257),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1257.INIT = 16'h8000;
LUT4 lut_inst_1258 (
  .F(lut_f_1258),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1258.INIT = 16'h8000;
LUT4 lut_inst_1259 (
  .F(lut_f_1259),
  .I0(lut_f_1256),
  .I1(lut_f_1257),
  .I2(lut_f_1258),
  .I3(gw_vcc)
);
defparam lut_inst_1259.INIT = 16'h8000;
LUT4 lut_inst_1260 (
  .F(lut_f_1260),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1260.INIT = 16'h8000;
LUT4 lut_inst_1261 (
  .F(lut_f_1261),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1261.INIT = 16'h8000;
LUT4 lut_inst_1262 (
  .F(lut_f_1262),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1262.INIT = 16'h8000;
LUT4 lut_inst_1263 (
  .F(lut_f_1263),
  .I0(lut_f_1260),
  .I1(lut_f_1261),
  .I2(lut_f_1262),
  .I3(gw_vcc)
);
defparam lut_inst_1263.INIT = 16'h8000;
LUT4 lut_inst_1264 (
  .F(lut_f_1264),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1264.INIT = 16'h8000;
LUT4 lut_inst_1265 (
  .F(lut_f_1265),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1265.INIT = 16'h8000;
LUT4 lut_inst_1266 (
  .F(lut_f_1266),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1266.INIT = 16'h8000;
LUT4 lut_inst_1267 (
  .F(lut_f_1267),
  .I0(lut_f_1264),
  .I1(lut_f_1265),
  .I2(lut_f_1266),
  .I3(gw_vcc)
);
defparam lut_inst_1267.INIT = 16'h8000;
LUT4 lut_inst_1268 (
  .F(lut_f_1268),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1268.INIT = 16'h8000;
LUT4 lut_inst_1269 (
  .F(lut_f_1269),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1269.INIT = 16'h8000;
LUT4 lut_inst_1270 (
  .F(lut_f_1270),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1270.INIT = 16'h8000;
LUT4 lut_inst_1271 (
  .F(lut_f_1271),
  .I0(lut_f_1268),
  .I1(lut_f_1269),
  .I2(lut_f_1270),
  .I3(gw_vcc)
);
defparam lut_inst_1271.INIT = 16'h8000;
LUT4 lut_inst_1272 (
  .F(lut_f_1272),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1272.INIT = 16'h8000;
LUT4 lut_inst_1273 (
  .F(lut_f_1273),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1273.INIT = 16'h8000;
LUT4 lut_inst_1274 (
  .F(lut_f_1274),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1274.INIT = 16'h8000;
LUT4 lut_inst_1275 (
  .F(lut_f_1275),
  .I0(lut_f_1272),
  .I1(lut_f_1273),
  .I2(lut_f_1274),
  .I3(gw_vcc)
);
defparam lut_inst_1275.INIT = 16'h8000;
LUT4 lut_inst_1276 (
  .F(lut_f_1276),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1276.INIT = 16'h8000;
LUT4 lut_inst_1277 (
  .F(lut_f_1277),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1277.INIT = 16'h8000;
LUT4 lut_inst_1278 (
  .F(lut_f_1278),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1278.INIT = 16'h8000;
LUT4 lut_inst_1279 (
  .F(lut_f_1279),
  .I0(lut_f_1276),
  .I1(lut_f_1277),
  .I2(lut_f_1278),
  .I3(gw_vcc)
);
defparam lut_inst_1279.INIT = 16'h8000;
LUT4 lut_inst_1280 (
  .F(lut_f_1280),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1280.INIT = 16'h8000;
LUT4 lut_inst_1281 (
  .F(lut_f_1281),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1281.INIT = 16'h8000;
LUT4 lut_inst_1282 (
  .F(lut_f_1282),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1282.INIT = 16'h8000;
LUT4 lut_inst_1283 (
  .F(lut_f_1283),
  .I0(lut_f_1280),
  .I1(lut_f_1281),
  .I2(lut_f_1282),
  .I3(gw_vcc)
);
defparam lut_inst_1283.INIT = 16'h8000;
LUT4 lut_inst_1284 (
  .F(lut_f_1284),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1284.INIT = 16'h8000;
LUT4 lut_inst_1285 (
  .F(lut_f_1285),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1285.INIT = 16'h8000;
LUT4 lut_inst_1286 (
  .F(lut_f_1286),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1286.INIT = 16'h8000;
LUT4 lut_inst_1287 (
  .F(lut_f_1287),
  .I0(lut_f_1284),
  .I1(lut_f_1285),
  .I2(lut_f_1286),
  .I3(gw_vcc)
);
defparam lut_inst_1287.INIT = 16'h8000;
LUT4 lut_inst_1288 (
  .F(lut_f_1288),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1288.INIT = 16'h8000;
LUT4 lut_inst_1289 (
  .F(lut_f_1289),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1289.INIT = 16'h8000;
LUT4 lut_inst_1290 (
  .F(lut_f_1290),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1290.INIT = 16'h8000;
LUT4 lut_inst_1291 (
  .F(lut_f_1291),
  .I0(lut_f_1288),
  .I1(lut_f_1289),
  .I2(lut_f_1290),
  .I3(gw_vcc)
);
defparam lut_inst_1291.INIT = 16'h8000;
LUT4 lut_inst_1292 (
  .F(lut_f_1292),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1292.INIT = 16'h8000;
LUT4 lut_inst_1293 (
  .F(lut_f_1293),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1293.INIT = 16'h8000;
LUT4 lut_inst_1294 (
  .F(lut_f_1294),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1294.INIT = 16'h8000;
LUT4 lut_inst_1295 (
  .F(lut_f_1295),
  .I0(lut_f_1292),
  .I1(lut_f_1293),
  .I2(lut_f_1294),
  .I3(gw_vcc)
);
defparam lut_inst_1295.INIT = 16'h8000;
LUT4 lut_inst_1296 (
  .F(lut_f_1296),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1296.INIT = 16'h8000;
LUT4 lut_inst_1297 (
  .F(lut_f_1297),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1297.INIT = 16'h8000;
LUT4 lut_inst_1298 (
  .F(lut_f_1298),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1298.INIT = 16'h8000;
LUT4 lut_inst_1299 (
  .F(lut_f_1299),
  .I0(lut_f_1296),
  .I1(lut_f_1297),
  .I2(lut_f_1298),
  .I3(gw_vcc)
);
defparam lut_inst_1299.INIT = 16'h8000;
LUT4 lut_inst_1300 (
  .F(lut_f_1300),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1300.INIT = 16'h8000;
LUT4 lut_inst_1301 (
  .F(lut_f_1301),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1301.INIT = 16'h8000;
LUT4 lut_inst_1302 (
  .F(lut_f_1302),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1302.INIT = 16'h8000;
LUT4 lut_inst_1303 (
  .F(lut_f_1303),
  .I0(lut_f_1300),
  .I1(lut_f_1301),
  .I2(lut_f_1302),
  .I3(gw_vcc)
);
defparam lut_inst_1303.INIT = 16'h8000;
LUT4 lut_inst_1304 (
  .F(lut_f_1304),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1304.INIT = 16'h8000;
LUT4 lut_inst_1305 (
  .F(lut_f_1305),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1305.INIT = 16'h8000;
LUT4 lut_inst_1306 (
  .F(lut_f_1306),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1306.INIT = 16'h8000;
LUT4 lut_inst_1307 (
  .F(lut_f_1307),
  .I0(lut_f_1304),
  .I1(lut_f_1305),
  .I2(lut_f_1306),
  .I3(gw_vcc)
);
defparam lut_inst_1307.INIT = 16'h8000;
LUT4 lut_inst_1308 (
  .F(lut_f_1308),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1308.INIT = 16'h8000;
LUT4 lut_inst_1309 (
  .F(lut_f_1309),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1309.INIT = 16'h8000;
LUT4 lut_inst_1310 (
  .F(lut_f_1310),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1310.INIT = 16'h8000;
LUT4 lut_inst_1311 (
  .F(lut_f_1311),
  .I0(lut_f_1308),
  .I1(lut_f_1309),
  .I2(lut_f_1310),
  .I3(gw_vcc)
);
defparam lut_inst_1311.INIT = 16'h8000;
LUT4 lut_inst_1312 (
  .F(lut_f_1312),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1312.INIT = 16'h8000;
LUT4 lut_inst_1313 (
  .F(lut_f_1313),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1313.INIT = 16'h8000;
LUT4 lut_inst_1314 (
  .F(lut_f_1314),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1314.INIT = 16'h8000;
LUT4 lut_inst_1315 (
  .F(lut_f_1315),
  .I0(lut_f_1312),
  .I1(lut_f_1313),
  .I2(lut_f_1314),
  .I3(gw_vcc)
);
defparam lut_inst_1315.INIT = 16'h8000;
LUT4 lut_inst_1316 (
  .F(lut_f_1316),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1316.INIT = 16'h8000;
LUT4 lut_inst_1317 (
  .F(lut_f_1317),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1317.INIT = 16'h8000;
LUT4 lut_inst_1318 (
  .F(lut_f_1318),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1318.INIT = 16'h8000;
LUT4 lut_inst_1319 (
  .F(lut_f_1319),
  .I0(lut_f_1316),
  .I1(lut_f_1317),
  .I2(lut_f_1318),
  .I3(gw_vcc)
);
defparam lut_inst_1319.INIT = 16'h8000;
LUT4 lut_inst_1320 (
  .F(lut_f_1320),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1320.INIT = 16'h8000;
LUT4 lut_inst_1321 (
  .F(lut_f_1321),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1321.INIT = 16'h8000;
LUT4 lut_inst_1322 (
  .F(lut_f_1322),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1322.INIT = 16'h8000;
LUT4 lut_inst_1323 (
  .F(lut_f_1323),
  .I0(lut_f_1320),
  .I1(lut_f_1321),
  .I2(lut_f_1322),
  .I3(gw_vcc)
);
defparam lut_inst_1323.INIT = 16'h8000;
LUT4 lut_inst_1324 (
  .F(lut_f_1324),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1324.INIT = 16'h8000;
LUT4 lut_inst_1325 (
  .F(lut_f_1325),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1325.INIT = 16'h8000;
LUT4 lut_inst_1326 (
  .F(lut_f_1326),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1326.INIT = 16'h8000;
LUT4 lut_inst_1327 (
  .F(lut_f_1327),
  .I0(lut_f_1324),
  .I1(lut_f_1325),
  .I2(lut_f_1326),
  .I3(gw_vcc)
);
defparam lut_inst_1327.INIT = 16'h8000;
LUT4 lut_inst_1328 (
  .F(lut_f_1328),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1328.INIT = 16'h8000;
LUT4 lut_inst_1329 (
  .F(lut_f_1329),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1329.INIT = 16'h8000;
LUT4 lut_inst_1330 (
  .F(lut_f_1330),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1330.INIT = 16'h8000;
LUT4 lut_inst_1331 (
  .F(lut_f_1331),
  .I0(lut_f_1328),
  .I1(lut_f_1329),
  .I2(lut_f_1330),
  .I3(gw_vcc)
);
defparam lut_inst_1331.INIT = 16'h8000;
LUT4 lut_inst_1332 (
  .F(lut_f_1332),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1332.INIT = 16'h8000;
LUT4 lut_inst_1333 (
  .F(lut_f_1333),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1333.INIT = 16'h8000;
LUT4 lut_inst_1334 (
  .F(lut_f_1334),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1334.INIT = 16'h8000;
LUT4 lut_inst_1335 (
  .F(lut_f_1335),
  .I0(lut_f_1332),
  .I1(lut_f_1333),
  .I2(lut_f_1334),
  .I3(gw_vcc)
);
defparam lut_inst_1335.INIT = 16'h8000;
LUT4 lut_inst_1336 (
  .F(lut_f_1336),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1336.INIT = 16'h8000;
LUT4 lut_inst_1337 (
  .F(lut_f_1337),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1337.INIT = 16'h8000;
LUT4 lut_inst_1338 (
  .F(lut_f_1338),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1338.INIT = 16'h8000;
LUT4 lut_inst_1339 (
  .F(lut_f_1339),
  .I0(lut_f_1336),
  .I1(lut_f_1337),
  .I2(lut_f_1338),
  .I3(gw_vcc)
);
defparam lut_inst_1339.INIT = 16'h8000;
LUT4 lut_inst_1340 (
  .F(lut_f_1340),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1340.INIT = 16'h8000;
LUT4 lut_inst_1341 (
  .F(lut_f_1341),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1341.INIT = 16'h8000;
LUT4 lut_inst_1342 (
  .F(lut_f_1342),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1342.INIT = 16'h8000;
LUT4 lut_inst_1343 (
  .F(lut_f_1343),
  .I0(lut_f_1340),
  .I1(lut_f_1341),
  .I2(lut_f_1342),
  .I3(gw_vcc)
);
defparam lut_inst_1343.INIT = 16'h8000;
LUT4 lut_inst_1344 (
  .F(lut_f_1344),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1344.INIT = 16'h8000;
LUT4 lut_inst_1345 (
  .F(lut_f_1345),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1345.INIT = 16'h8000;
LUT4 lut_inst_1346 (
  .F(lut_f_1346),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1346.INIT = 16'h8000;
LUT4 lut_inst_1347 (
  .F(lut_f_1347),
  .I0(lut_f_1344),
  .I1(lut_f_1345),
  .I2(lut_f_1346),
  .I3(gw_vcc)
);
defparam lut_inst_1347.INIT = 16'h8000;
LUT4 lut_inst_1348 (
  .F(lut_f_1348),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1348.INIT = 16'h8000;
LUT4 lut_inst_1349 (
  .F(lut_f_1349),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1349.INIT = 16'h8000;
LUT4 lut_inst_1350 (
  .F(lut_f_1350),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1350.INIT = 16'h8000;
LUT4 lut_inst_1351 (
  .F(lut_f_1351),
  .I0(lut_f_1348),
  .I1(lut_f_1349),
  .I2(lut_f_1350),
  .I3(gw_vcc)
);
defparam lut_inst_1351.INIT = 16'h8000;
LUT4 lut_inst_1352 (
  .F(lut_f_1352),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1352.INIT = 16'h8000;
LUT4 lut_inst_1353 (
  .F(lut_f_1353),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1353.INIT = 16'h8000;
LUT4 lut_inst_1354 (
  .F(lut_f_1354),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1354.INIT = 16'h8000;
LUT4 lut_inst_1355 (
  .F(lut_f_1355),
  .I0(lut_f_1352),
  .I1(lut_f_1353),
  .I2(lut_f_1354),
  .I3(gw_vcc)
);
defparam lut_inst_1355.INIT = 16'h8000;
LUT4 lut_inst_1356 (
  .F(lut_f_1356),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1356.INIT = 16'h8000;
LUT4 lut_inst_1357 (
  .F(lut_f_1357),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1357.INIT = 16'h8000;
LUT4 lut_inst_1358 (
  .F(lut_f_1358),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1358.INIT = 16'h8000;
LUT4 lut_inst_1359 (
  .F(lut_f_1359),
  .I0(lut_f_1356),
  .I1(lut_f_1357),
  .I2(lut_f_1358),
  .I3(gw_vcc)
);
defparam lut_inst_1359.INIT = 16'h8000;
LUT4 lut_inst_1360 (
  .F(lut_f_1360),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1360.INIT = 16'h8000;
LUT4 lut_inst_1361 (
  .F(lut_f_1361),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1361.INIT = 16'h8000;
LUT4 lut_inst_1362 (
  .F(lut_f_1362),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1362.INIT = 16'h8000;
LUT4 lut_inst_1363 (
  .F(lut_f_1363),
  .I0(lut_f_1360),
  .I1(lut_f_1361),
  .I2(lut_f_1362),
  .I3(gw_vcc)
);
defparam lut_inst_1363.INIT = 16'h8000;
LUT4 lut_inst_1364 (
  .F(lut_f_1364),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1364.INIT = 16'h8000;
LUT4 lut_inst_1365 (
  .F(lut_f_1365),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1365.INIT = 16'h8000;
LUT4 lut_inst_1366 (
  .F(lut_f_1366),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1366.INIT = 16'h8000;
LUT4 lut_inst_1367 (
  .F(lut_f_1367),
  .I0(lut_f_1364),
  .I1(lut_f_1365),
  .I2(lut_f_1366),
  .I3(gw_vcc)
);
defparam lut_inst_1367.INIT = 16'h8000;
LUT4 lut_inst_1368 (
  .F(lut_f_1368),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1368.INIT = 16'h8000;
LUT4 lut_inst_1369 (
  .F(lut_f_1369),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1369.INIT = 16'h8000;
LUT4 lut_inst_1370 (
  .F(lut_f_1370),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1370.INIT = 16'h8000;
LUT4 lut_inst_1371 (
  .F(lut_f_1371),
  .I0(lut_f_1368),
  .I1(lut_f_1369),
  .I2(lut_f_1370),
  .I3(gw_vcc)
);
defparam lut_inst_1371.INIT = 16'h8000;
LUT4 lut_inst_1372 (
  .F(lut_f_1372),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1372.INIT = 16'h8000;
LUT4 lut_inst_1373 (
  .F(lut_f_1373),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1373.INIT = 16'h8000;
LUT4 lut_inst_1374 (
  .F(lut_f_1374),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1374.INIT = 16'h8000;
LUT4 lut_inst_1375 (
  .F(lut_f_1375),
  .I0(lut_f_1372),
  .I1(lut_f_1373),
  .I2(lut_f_1374),
  .I3(gw_vcc)
);
defparam lut_inst_1375.INIT = 16'h8000;
LUT4 lut_inst_1376 (
  .F(lut_f_1376),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1376.INIT = 16'h8000;
LUT4 lut_inst_1377 (
  .F(lut_f_1377),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1377.INIT = 16'h8000;
LUT4 lut_inst_1378 (
  .F(lut_f_1378),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1378.INIT = 16'h8000;
LUT4 lut_inst_1379 (
  .F(lut_f_1379),
  .I0(lut_f_1376),
  .I1(lut_f_1377),
  .I2(lut_f_1378),
  .I3(gw_vcc)
);
defparam lut_inst_1379.INIT = 16'h8000;
LUT4 lut_inst_1380 (
  .F(lut_f_1380),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1380.INIT = 16'h8000;
LUT4 lut_inst_1381 (
  .F(lut_f_1381),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1381.INIT = 16'h8000;
LUT4 lut_inst_1382 (
  .F(lut_f_1382),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1382.INIT = 16'h8000;
LUT4 lut_inst_1383 (
  .F(lut_f_1383),
  .I0(lut_f_1380),
  .I1(lut_f_1381),
  .I2(lut_f_1382),
  .I3(gw_vcc)
);
defparam lut_inst_1383.INIT = 16'h8000;
LUT4 lut_inst_1384 (
  .F(lut_f_1384),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1384.INIT = 16'h8000;
LUT4 lut_inst_1385 (
  .F(lut_f_1385),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1385.INIT = 16'h8000;
LUT4 lut_inst_1386 (
  .F(lut_f_1386),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1386.INIT = 16'h8000;
LUT4 lut_inst_1387 (
  .F(lut_f_1387),
  .I0(lut_f_1384),
  .I1(lut_f_1385),
  .I2(lut_f_1386),
  .I3(gw_vcc)
);
defparam lut_inst_1387.INIT = 16'h8000;
LUT4 lut_inst_1388 (
  .F(lut_f_1388),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1388.INIT = 16'h8000;
LUT4 lut_inst_1389 (
  .F(lut_f_1389),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1389.INIT = 16'h8000;
LUT4 lut_inst_1390 (
  .F(lut_f_1390),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1390.INIT = 16'h8000;
LUT4 lut_inst_1391 (
  .F(lut_f_1391),
  .I0(lut_f_1388),
  .I1(lut_f_1389),
  .I2(lut_f_1390),
  .I3(gw_vcc)
);
defparam lut_inst_1391.INIT = 16'h8000;
LUT4 lut_inst_1392 (
  .F(lut_f_1392),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1392.INIT = 16'h8000;
LUT4 lut_inst_1393 (
  .F(lut_f_1393),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1393.INIT = 16'h8000;
LUT4 lut_inst_1394 (
  .F(lut_f_1394),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1394.INIT = 16'h8000;
LUT4 lut_inst_1395 (
  .F(lut_f_1395),
  .I0(lut_f_1392),
  .I1(lut_f_1393),
  .I2(lut_f_1394),
  .I3(gw_vcc)
);
defparam lut_inst_1395.INIT = 16'h8000;
LUT4 lut_inst_1396 (
  .F(lut_f_1396),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1396.INIT = 16'h8000;
LUT4 lut_inst_1397 (
  .F(lut_f_1397),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1397.INIT = 16'h8000;
LUT4 lut_inst_1398 (
  .F(lut_f_1398),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1398.INIT = 16'h8000;
LUT4 lut_inst_1399 (
  .F(lut_f_1399),
  .I0(lut_f_1396),
  .I1(lut_f_1397),
  .I2(lut_f_1398),
  .I3(gw_vcc)
);
defparam lut_inst_1399.INIT = 16'h8000;
LUT4 lut_inst_1400 (
  .F(lut_f_1400),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1400.INIT = 16'h8000;
LUT4 lut_inst_1401 (
  .F(lut_f_1401),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1401.INIT = 16'h8000;
LUT4 lut_inst_1402 (
  .F(lut_f_1402),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1402.INIT = 16'h8000;
LUT4 lut_inst_1403 (
  .F(lut_f_1403),
  .I0(lut_f_1400),
  .I1(lut_f_1401),
  .I2(lut_f_1402),
  .I3(gw_vcc)
);
defparam lut_inst_1403.INIT = 16'h8000;
LUT4 lut_inst_1404 (
  .F(lut_f_1404),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1404.INIT = 16'h8000;
LUT4 lut_inst_1405 (
  .F(lut_f_1405),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1405.INIT = 16'h8000;
LUT4 lut_inst_1406 (
  .F(lut_f_1406),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1406.INIT = 16'h8000;
LUT4 lut_inst_1407 (
  .F(lut_f_1407),
  .I0(lut_f_1404),
  .I1(lut_f_1405),
  .I2(lut_f_1406),
  .I3(gw_vcc)
);
defparam lut_inst_1407.INIT = 16'h8000;
LUT4 lut_inst_1408 (
  .F(lut_f_1408),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1408.INIT = 16'h8000;
LUT4 lut_inst_1409 (
  .F(lut_f_1409),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1409.INIT = 16'h8000;
LUT4 lut_inst_1410 (
  .F(lut_f_1410),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1410.INIT = 16'h8000;
LUT4 lut_inst_1411 (
  .F(lut_f_1411),
  .I0(lut_f_1408),
  .I1(lut_f_1409),
  .I2(lut_f_1410),
  .I3(gw_vcc)
);
defparam lut_inst_1411.INIT = 16'h8000;
LUT4 lut_inst_1412 (
  .F(lut_f_1412),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1412.INIT = 16'h8000;
LUT4 lut_inst_1413 (
  .F(lut_f_1413),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1413.INIT = 16'h8000;
LUT4 lut_inst_1414 (
  .F(lut_f_1414),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1414.INIT = 16'h8000;
LUT4 lut_inst_1415 (
  .F(lut_f_1415),
  .I0(lut_f_1412),
  .I1(lut_f_1413),
  .I2(lut_f_1414),
  .I3(gw_vcc)
);
defparam lut_inst_1415.INIT = 16'h8000;
LUT4 lut_inst_1416 (
  .F(lut_f_1416),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1416.INIT = 16'h8000;
LUT4 lut_inst_1417 (
  .F(lut_f_1417),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1417.INIT = 16'h8000;
LUT4 lut_inst_1418 (
  .F(lut_f_1418),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1418.INIT = 16'h8000;
LUT4 lut_inst_1419 (
  .F(lut_f_1419),
  .I0(lut_f_1416),
  .I1(lut_f_1417),
  .I2(lut_f_1418),
  .I3(gw_vcc)
);
defparam lut_inst_1419.INIT = 16'h8000;
LUT4 lut_inst_1420 (
  .F(lut_f_1420),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1420.INIT = 16'h8000;
LUT4 lut_inst_1421 (
  .F(lut_f_1421),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1421.INIT = 16'h8000;
LUT4 lut_inst_1422 (
  .F(lut_f_1422),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1422.INIT = 16'h8000;
LUT4 lut_inst_1423 (
  .F(lut_f_1423),
  .I0(lut_f_1420),
  .I1(lut_f_1421),
  .I2(lut_f_1422),
  .I3(gw_vcc)
);
defparam lut_inst_1423.INIT = 16'h8000;
LUT4 lut_inst_1424 (
  .F(lut_f_1424),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1424.INIT = 16'h8000;
LUT4 lut_inst_1425 (
  .F(lut_f_1425),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1425.INIT = 16'h8000;
LUT4 lut_inst_1426 (
  .F(lut_f_1426),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1426.INIT = 16'h8000;
LUT4 lut_inst_1427 (
  .F(lut_f_1427),
  .I0(lut_f_1424),
  .I1(lut_f_1425),
  .I2(lut_f_1426),
  .I3(gw_vcc)
);
defparam lut_inst_1427.INIT = 16'h8000;
LUT4 lut_inst_1428 (
  .F(lut_f_1428),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1428.INIT = 16'h8000;
LUT4 lut_inst_1429 (
  .F(lut_f_1429),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1429.INIT = 16'h8000;
LUT4 lut_inst_1430 (
  .F(lut_f_1430),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1430.INIT = 16'h8000;
LUT4 lut_inst_1431 (
  .F(lut_f_1431),
  .I0(lut_f_1428),
  .I1(lut_f_1429),
  .I2(lut_f_1430),
  .I3(gw_vcc)
);
defparam lut_inst_1431.INIT = 16'h8000;
LUT4 lut_inst_1432 (
  .F(lut_f_1432),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1432.INIT = 16'h8000;
LUT4 lut_inst_1433 (
  .F(lut_f_1433),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1433.INIT = 16'h8000;
LUT4 lut_inst_1434 (
  .F(lut_f_1434),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1434.INIT = 16'h8000;
LUT4 lut_inst_1435 (
  .F(lut_f_1435),
  .I0(lut_f_1432),
  .I1(lut_f_1433),
  .I2(lut_f_1434),
  .I3(gw_vcc)
);
defparam lut_inst_1435.INIT = 16'h8000;
LUT4 lut_inst_1436 (
  .F(lut_f_1436),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1436.INIT = 16'h8000;
LUT4 lut_inst_1437 (
  .F(lut_f_1437),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1437.INIT = 16'h8000;
LUT4 lut_inst_1438 (
  .F(lut_f_1438),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1438.INIT = 16'h8000;
LUT4 lut_inst_1439 (
  .F(lut_f_1439),
  .I0(lut_f_1436),
  .I1(lut_f_1437),
  .I2(lut_f_1438),
  .I3(gw_vcc)
);
defparam lut_inst_1439.INIT = 16'h8000;
LUT4 lut_inst_1440 (
  .F(lut_f_1440),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1440.INIT = 16'h8000;
LUT4 lut_inst_1441 (
  .F(lut_f_1441),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1441.INIT = 16'h8000;
LUT4 lut_inst_1442 (
  .F(lut_f_1442),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1442.INIT = 16'h8000;
LUT4 lut_inst_1443 (
  .F(lut_f_1443),
  .I0(lut_f_1440),
  .I1(lut_f_1441),
  .I2(lut_f_1442),
  .I3(gw_vcc)
);
defparam lut_inst_1443.INIT = 16'h8000;
LUT4 lut_inst_1444 (
  .F(lut_f_1444),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1444.INIT = 16'h8000;
LUT4 lut_inst_1445 (
  .F(lut_f_1445),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1445.INIT = 16'h8000;
LUT4 lut_inst_1446 (
  .F(lut_f_1446),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1446.INIT = 16'h8000;
LUT4 lut_inst_1447 (
  .F(lut_f_1447),
  .I0(lut_f_1444),
  .I1(lut_f_1445),
  .I2(lut_f_1446),
  .I3(gw_vcc)
);
defparam lut_inst_1447.INIT = 16'h8000;
LUT4 lut_inst_1448 (
  .F(lut_f_1448),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1448.INIT = 16'h8000;
LUT4 lut_inst_1449 (
  .F(lut_f_1449),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1449.INIT = 16'h8000;
LUT4 lut_inst_1450 (
  .F(lut_f_1450),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1450.INIT = 16'h8000;
LUT4 lut_inst_1451 (
  .F(lut_f_1451),
  .I0(lut_f_1448),
  .I1(lut_f_1449),
  .I2(lut_f_1450),
  .I3(gw_vcc)
);
defparam lut_inst_1451.INIT = 16'h8000;
LUT4 lut_inst_1452 (
  .F(lut_f_1452),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1452.INIT = 16'h8000;
LUT4 lut_inst_1453 (
  .F(lut_f_1453),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1453.INIT = 16'h8000;
LUT4 lut_inst_1454 (
  .F(lut_f_1454),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1454.INIT = 16'h8000;
LUT4 lut_inst_1455 (
  .F(lut_f_1455),
  .I0(lut_f_1452),
  .I1(lut_f_1453),
  .I2(lut_f_1454),
  .I3(gw_vcc)
);
defparam lut_inst_1455.INIT = 16'h8000;
LUT4 lut_inst_1456 (
  .F(lut_f_1456),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1456.INIT = 16'h8000;
LUT4 lut_inst_1457 (
  .F(lut_f_1457),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1457.INIT = 16'h8000;
LUT4 lut_inst_1458 (
  .F(lut_f_1458),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1458.INIT = 16'h8000;
LUT4 lut_inst_1459 (
  .F(lut_f_1459),
  .I0(lut_f_1456),
  .I1(lut_f_1457),
  .I2(lut_f_1458),
  .I3(gw_vcc)
);
defparam lut_inst_1459.INIT = 16'h8000;
LUT4 lut_inst_1460 (
  .F(lut_f_1460),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1460.INIT = 16'h8000;
LUT4 lut_inst_1461 (
  .F(lut_f_1461),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1461.INIT = 16'h8000;
LUT4 lut_inst_1462 (
  .F(lut_f_1462),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1462.INIT = 16'h8000;
LUT4 lut_inst_1463 (
  .F(lut_f_1463),
  .I0(lut_f_1460),
  .I1(lut_f_1461),
  .I2(lut_f_1462),
  .I3(gw_vcc)
);
defparam lut_inst_1463.INIT = 16'h8000;
LUT4 lut_inst_1464 (
  .F(lut_f_1464),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1464.INIT = 16'h8000;
LUT4 lut_inst_1465 (
  .F(lut_f_1465),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1465.INIT = 16'h8000;
LUT4 lut_inst_1466 (
  .F(lut_f_1466),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1466.INIT = 16'h8000;
LUT4 lut_inst_1467 (
  .F(lut_f_1467),
  .I0(lut_f_1464),
  .I1(lut_f_1465),
  .I2(lut_f_1466),
  .I3(gw_vcc)
);
defparam lut_inst_1467.INIT = 16'h8000;
LUT4 lut_inst_1468 (
  .F(lut_f_1468),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1468.INIT = 16'h8000;
LUT4 lut_inst_1469 (
  .F(lut_f_1469),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1469.INIT = 16'h8000;
LUT4 lut_inst_1470 (
  .F(lut_f_1470),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1470.INIT = 16'h8000;
LUT4 lut_inst_1471 (
  .F(lut_f_1471),
  .I0(lut_f_1468),
  .I1(lut_f_1469),
  .I2(lut_f_1470),
  .I3(gw_vcc)
);
defparam lut_inst_1471.INIT = 16'h8000;
LUT4 lut_inst_1472 (
  .F(lut_f_1472),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1472.INIT = 16'h8000;
LUT4 lut_inst_1473 (
  .F(lut_f_1473),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1473.INIT = 16'h8000;
LUT4 lut_inst_1474 (
  .F(lut_f_1474),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1474.INIT = 16'h8000;
LUT4 lut_inst_1475 (
  .F(lut_f_1475),
  .I0(lut_f_1472),
  .I1(lut_f_1473),
  .I2(lut_f_1474),
  .I3(gw_vcc)
);
defparam lut_inst_1475.INIT = 16'h8000;
LUT4 lut_inst_1476 (
  .F(lut_f_1476),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1476.INIT = 16'h8000;
LUT4 lut_inst_1477 (
  .F(lut_f_1477),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1477.INIT = 16'h8000;
LUT4 lut_inst_1478 (
  .F(lut_f_1478),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1478.INIT = 16'h8000;
LUT4 lut_inst_1479 (
  .F(lut_f_1479),
  .I0(lut_f_1476),
  .I1(lut_f_1477),
  .I2(lut_f_1478),
  .I3(gw_vcc)
);
defparam lut_inst_1479.INIT = 16'h8000;
LUT4 lut_inst_1480 (
  .F(lut_f_1480),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1480.INIT = 16'h8000;
LUT4 lut_inst_1481 (
  .F(lut_f_1481),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1481.INIT = 16'h8000;
LUT4 lut_inst_1482 (
  .F(lut_f_1482),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1482.INIT = 16'h8000;
LUT4 lut_inst_1483 (
  .F(lut_f_1483),
  .I0(lut_f_1480),
  .I1(lut_f_1481),
  .I2(lut_f_1482),
  .I3(gw_vcc)
);
defparam lut_inst_1483.INIT = 16'h8000;
LUT4 lut_inst_1484 (
  .F(lut_f_1484),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1484.INIT = 16'h8000;
LUT4 lut_inst_1485 (
  .F(lut_f_1485),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1485.INIT = 16'h8000;
LUT4 lut_inst_1486 (
  .F(lut_f_1486),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1486.INIT = 16'h8000;
LUT4 lut_inst_1487 (
  .F(lut_f_1487),
  .I0(lut_f_1484),
  .I1(lut_f_1485),
  .I2(lut_f_1486),
  .I3(gw_vcc)
);
defparam lut_inst_1487.INIT = 16'h8000;
LUT4 lut_inst_1488 (
  .F(lut_f_1488),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1488.INIT = 16'h8000;
LUT4 lut_inst_1489 (
  .F(lut_f_1489),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1489.INIT = 16'h8000;
LUT4 lut_inst_1490 (
  .F(lut_f_1490),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1490.INIT = 16'h8000;
LUT4 lut_inst_1491 (
  .F(lut_f_1491),
  .I0(lut_f_1488),
  .I1(lut_f_1489),
  .I2(lut_f_1490),
  .I3(gw_vcc)
);
defparam lut_inst_1491.INIT = 16'h8000;
LUT4 lut_inst_1492 (
  .F(lut_f_1492),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1492.INIT = 16'h8000;
LUT4 lut_inst_1493 (
  .F(lut_f_1493),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1493.INIT = 16'h8000;
LUT4 lut_inst_1494 (
  .F(lut_f_1494),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1494.INIT = 16'h8000;
LUT4 lut_inst_1495 (
  .F(lut_f_1495),
  .I0(lut_f_1492),
  .I1(lut_f_1493),
  .I2(lut_f_1494),
  .I3(gw_vcc)
);
defparam lut_inst_1495.INIT = 16'h8000;
LUT4 lut_inst_1496 (
  .F(lut_f_1496),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1496.INIT = 16'h8000;
LUT4 lut_inst_1497 (
  .F(lut_f_1497),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1497.INIT = 16'h8000;
LUT4 lut_inst_1498 (
  .F(lut_f_1498),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1498.INIT = 16'h8000;
LUT4 lut_inst_1499 (
  .F(lut_f_1499),
  .I0(lut_f_1496),
  .I1(lut_f_1497),
  .I2(lut_f_1498),
  .I3(gw_vcc)
);
defparam lut_inst_1499.INIT = 16'h8000;
LUT4 lut_inst_1500 (
  .F(lut_f_1500),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1500.INIT = 16'h8000;
LUT4 lut_inst_1501 (
  .F(lut_f_1501),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1501.INIT = 16'h8000;
LUT4 lut_inst_1502 (
  .F(lut_f_1502),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1502.INIT = 16'h8000;
LUT4 lut_inst_1503 (
  .F(lut_f_1503),
  .I0(lut_f_1500),
  .I1(lut_f_1501),
  .I2(lut_f_1502),
  .I3(gw_vcc)
);
defparam lut_inst_1503.INIT = 16'h8000;
LUT4 lut_inst_1504 (
  .F(lut_f_1504),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1504.INIT = 16'h8000;
LUT4 lut_inst_1505 (
  .F(lut_f_1505),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1505.INIT = 16'h8000;
LUT4 lut_inst_1506 (
  .F(lut_f_1506),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1506.INIT = 16'h8000;
LUT4 lut_inst_1507 (
  .F(lut_f_1507),
  .I0(lut_f_1504),
  .I1(lut_f_1505),
  .I2(lut_f_1506),
  .I3(gw_vcc)
);
defparam lut_inst_1507.INIT = 16'h8000;
LUT4 lut_inst_1508 (
  .F(lut_f_1508),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1508.INIT = 16'h8000;
LUT4 lut_inst_1509 (
  .F(lut_f_1509),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1509.INIT = 16'h8000;
LUT4 lut_inst_1510 (
  .F(lut_f_1510),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1510.INIT = 16'h8000;
LUT4 lut_inst_1511 (
  .F(lut_f_1511),
  .I0(lut_f_1508),
  .I1(lut_f_1509),
  .I2(lut_f_1510),
  .I3(gw_vcc)
);
defparam lut_inst_1511.INIT = 16'h8000;
LUT4 lut_inst_1512 (
  .F(lut_f_1512),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1512.INIT = 16'h8000;
LUT4 lut_inst_1513 (
  .F(lut_f_1513),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1513.INIT = 16'h8000;
LUT4 lut_inst_1514 (
  .F(lut_f_1514),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1514.INIT = 16'h8000;
LUT4 lut_inst_1515 (
  .F(lut_f_1515),
  .I0(lut_f_1512),
  .I1(lut_f_1513),
  .I2(lut_f_1514),
  .I3(gw_vcc)
);
defparam lut_inst_1515.INIT = 16'h8000;
LUT4 lut_inst_1516 (
  .F(lut_f_1516),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1516.INIT = 16'h8000;
LUT4 lut_inst_1517 (
  .F(lut_f_1517),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1517.INIT = 16'h8000;
LUT4 lut_inst_1518 (
  .F(lut_f_1518),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1518.INIT = 16'h8000;
LUT4 lut_inst_1519 (
  .F(lut_f_1519),
  .I0(lut_f_1516),
  .I1(lut_f_1517),
  .I2(lut_f_1518),
  .I3(gw_vcc)
);
defparam lut_inst_1519.INIT = 16'h8000;
LUT4 lut_inst_1520 (
  .F(lut_f_1520),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1520.INIT = 16'h8000;
LUT4 lut_inst_1521 (
  .F(lut_f_1521),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1521.INIT = 16'h8000;
LUT4 lut_inst_1522 (
  .F(lut_f_1522),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1522.INIT = 16'h8000;
LUT4 lut_inst_1523 (
  .F(lut_f_1523),
  .I0(lut_f_1520),
  .I1(lut_f_1521),
  .I2(lut_f_1522),
  .I3(gw_vcc)
);
defparam lut_inst_1523.INIT = 16'h8000;
LUT4 lut_inst_1524 (
  .F(lut_f_1524),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1524.INIT = 16'h8000;
LUT4 lut_inst_1525 (
  .F(lut_f_1525),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1525.INIT = 16'h8000;
LUT4 lut_inst_1526 (
  .F(lut_f_1526),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1526.INIT = 16'h8000;
LUT4 lut_inst_1527 (
  .F(lut_f_1527),
  .I0(lut_f_1524),
  .I1(lut_f_1525),
  .I2(lut_f_1526),
  .I3(gw_vcc)
);
defparam lut_inst_1527.INIT = 16'h8000;
LUT4 lut_inst_1528 (
  .F(lut_f_1528),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1528.INIT = 16'h8000;
LUT4 lut_inst_1529 (
  .F(lut_f_1529),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1529.INIT = 16'h8000;
LUT4 lut_inst_1530 (
  .F(lut_f_1530),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1530.INIT = 16'h8000;
LUT4 lut_inst_1531 (
  .F(lut_f_1531),
  .I0(lut_f_1528),
  .I1(lut_f_1529),
  .I2(lut_f_1530),
  .I3(gw_vcc)
);
defparam lut_inst_1531.INIT = 16'h8000;
LUT4 lut_inst_1532 (
  .F(lut_f_1532),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1532.INIT = 16'h8000;
LUT4 lut_inst_1533 (
  .F(lut_f_1533),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1533.INIT = 16'h8000;
LUT4 lut_inst_1534 (
  .F(lut_f_1534),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1534.INIT = 16'h8000;
LUT4 lut_inst_1535 (
  .F(lut_f_1535),
  .I0(lut_f_1532),
  .I1(lut_f_1533),
  .I2(lut_f_1534),
  .I3(gw_vcc)
);
defparam lut_inst_1535.INIT = 16'h8000;
LUT4 lut_inst_1536 (
  .F(lut_f_1536),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1536.INIT = 16'h8000;
LUT4 lut_inst_1537 (
  .F(lut_f_1537),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1537.INIT = 16'h8000;
LUT4 lut_inst_1538 (
  .F(lut_f_1538),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1538.INIT = 16'h8000;
LUT4 lut_inst_1539 (
  .F(lut_f_1539),
  .I0(lut_f_1536),
  .I1(lut_f_1537),
  .I2(lut_f_1538),
  .I3(gw_vcc)
);
defparam lut_inst_1539.INIT = 16'h8000;
LUT4 lut_inst_1540 (
  .F(lut_f_1540),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1540.INIT = 16'h8000;
LUT4 lut_inst_1541 (
  .F(lut_f_1541),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1541.INIT = 16'h8000;
LUT4 lut_inst_1542 (
  .F(lut_f_1542),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1542.INIT = 16'h8000;
LUT4 lut_inst_1543 (
  .F(lut_f_1543),
  .I0(lut_f_1540),
  .I1(lut_f_1541),
  .I2(lut_f_1542),
  .I3(gw_vcc)
);
defparam lut_inst_1543.INIT = 16'h8000;
LUT4 lut_inst_1544 (
  .F(lut_f_1544),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1544.INIT = 16'h8000;
LUT4 lut_inst_1545 (
  .F(lut_f_1545),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1545.INIT = 16'h8000;
LUT4 lut_inst_1546 (
  .F(lut_f_1546),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1546.INIT = 16'h8000;
LUT4 lut_inst_1547 (
  .F(lut_f_1547),
  .I0(lut_f_1544),
  .I1(lut_f_1545),
  .I2(lut_f_1546),
  .I3(gw_vcc)
);
defparam lut_inst_1547.INIT = 16'h8000;
LUT4 lut_inst_1548 (
  .F(lut_f_1548),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1548.INIT = 16'h8000;
LUT4 lut_inst_1549 (
  .F(lut_f_1549),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1549.INIT = 16'h8000;
LUT4 lut_inst_1550 (
  .F(lut_f_1550),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1550.INIT = 16'h8000;
LUT4 lut_inst_1551 (
  .F(lut_f_1551),
  .I0(lut_f_1548),
  .I1(lut_f_1549),
  .I2(lut_f_1550),
  .I3(gw_vcc)
);
defparam lut_inst_1551.INIT = 16'h8000;
LUT4 lut_inst_1552 (
  .F(lut_f_1552),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1552.INIT = 16'h8000;
LUT4 lut_inst_1553 (
  .F(lut_f_1553),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1553.INIT = 16'h8000;
LUT4 lut_inst_1554 (
  .F(lut_f_1554),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1554.INIT = 16'h8000;
LUT4 lut_inst_1555 (
  .F(lut_f_1555),
  .I0(lut_f_1552),
  .I1(lut_f_1553),
  .I2(lut_f_1554),
  .I3(gw_vcc)
);
defparam lut_inst_1555.INIT = 16'h8000;
LUT4 lut_inst_1556 (
  .F(lut_f_1556),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1556.INIT = 16'h8000;
LUT4 lut_inst_1557 (
  .F(lut_f_1557),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1557.INIT = 16'h8000;
LUT4 lut_inst_1558 (
  .F(lut_f_1558),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1558.INIT = 16'h8000;
LUT4 lut_inst_1559 (
  .F(lut_f_1559),
  .I0(lut_f_1556),
  .I1(lut_f_1557),
  .I2(lut_f_1558),
  .I3(gw_vcc)
);
defparam lut_inst_1559.INIT = 16'h8000;
LUT4 lut_inst_1560 (
  .F(lut_f_1560),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1560.INIT = 16'h8000;
LUT4 lut_inst_1561 (
  .F(lut_f_1561),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1561.INIT = 16'h8000;
LUT4 lut_inst_1562 (
  .F(lut_f_1562),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1562.INIT = 16'h8000;
LUT4 lut_inst_1563 (
  .F(lut_f_1563),
  .I0(lut_f_1560),
  .I1(lut_f_1561),
  .I2(lut_f_1562),
  .I3(gw_vcc)
);
defparam lut_inst_1563.INIT = 16'h8000;
LUT4 lut_inst_1564 (
  .F(lut_f_1564),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1564.INIT = 16'h8000;
LUT4 lut_inst_1565 (
  .F(lut_f_1565),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1565.INIT = 16'h8000;
LUT4 lut_inst_1566 (
  .F(lut_f_1566),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1566.INIT = 16'h8000;
LUT4 lut_inst_1567 (
  .F(lut_f_1567),
  .I0(lut_f_1564),
  .I1(lut_f_1565),
  .I2(lut_f_1566),
  .I3(gw_vcc)
);
defparam lut_inst_1567.INIT = 16'h8000;
LUT4 lut_inst_1568 (
  .F(lut_f_1568),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1568.INIT = 16'h8000;
LUT4 lut_inst_1569 (
  .F(lut_f_1569),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1569.INIT = 16'h8000;
LUT4 lut_inst_1570 (
  .F(lut_f_1570),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1570.INIT = 16'h8000;
LUT4 lut_inst_1571 (
  .F(lut_f_1571),
  .I0(lut_f_1568),
  .I1(lut_f_1569),
  .I2(lut_f_1570),
  .I3(gw_vcc)
);
defparam lut_inst_1571.INIT = 16'h8000;
LUT4 lut_inst_1572 (
  .F(lut_f_1572),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1572.INIT = 16'h8000;
LUT4 lut_inst_1573 (
  .F(lut_f_1573),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1573.INIT = 16'h8000;
LUT4 lut_inst_1574 (
  .F(lut_f_1574),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1574.INIT = 16'h8000;
LUT4 lut_inst_1575 (
  .F(lut_f_1575),
  .I0(lut_f_1572),
  .I1(lut_f_1573),
  .I2(lut_f_1574),
  .I3(gw_vcc)
);
defparam lut_inst_1575.INIT = 16'h8000;
LUT4 lut_inst_1576 (
  .F(lut_f_1576),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1576.INIT = 16'h8000;
LUT4 lut_inst_1577 (
  .F(lut_f_1577),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1577.INIT = 16'h8000;
LUT4 lut_inst_1578 (
  .F(lut_f_1578),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1578.INIT = 16'h8000;
LUT4 lut_inst_1579 (
  .F(lut_f_1579),
  .I0(lut_f_1576),
  .I1(lut_f_1577),
  .I2(lut_f_1578),
  .I3(gw_vcc)
);
defparam lut_inst_1579.INIT = 16'h8000;
LUT4 lut_inst_1580 (
  .F(lut_f_1580),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1580.INIT = 16'h8000;
LUT4 lut_inst_1581 (
  .F(lut_f_1581),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1581.INIT = 16'h8000;
LUT4 lut_inst_1582 (
  .F(lut_f_1582),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1582.INIT = 16'h8000;
LUT4 lut_inst_1583 (
  .F(lut_f_1583),
  .I0(lut_f_1580),
  .I1(lut_f_1581),
  .I2(lut_f_1582),
  .I3(gw_vcc)
);
defparam lut_inst_1583.INIT = 16'h8000;
LUT4 lut_inst_1584 (
  .F(lut_f_1584),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1584.INIT = 16'h8000;
LUT4 lut_inst_1585 (
  .F(lut_f_1585),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1585.INIT = 16'h8000;
LUT4 lut_inst_1586 (
  .F(lut_f_1586),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1586.INIT = 16'h8000;
LUT4 lut_inst_1587 (
  .F(lut_f_1587),
  .I0(lut_f_1584),
  .I1(lut_f_1585),
  .I2(lut_f_1586),
  .I3(gw_vcc)
);
defparam lut_inst_1587.INIT = 16'h8000;
LUT4 lut_inst_1588 (
  .F(lut_f_1588),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1588.INIT = 16'h8000;
LUT4 lut_inst_1589 (
  .F(lut_f_1589),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1589.INIT = 16'h8000;
LUT4 lut_inst_1590 (
  .F(lut_f_1590),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1590.INIT = 16'h8000;
LUT4 lut_inst_1591 (
  .F(lut_f_1591),
  .I0(lut_f_1588),
  .I1(lut_f_1589),
  .I2(lut_f_1590),
  .I3(gw_vcc)
);
defparam lut_inst_1591.INIT = 16'h8000;
LUT4 lut_inst_1592 (
  .F(lut_f_1592),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1592.INIT = 16'h8000;
LUT4 lut_inst_1593 (
  .F(lut_f_1593),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1593.INIT = 16'h8000;
LUT4 lut_inst_1594 (
  .F(lut_f_1594),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1594.INIT = 16'h8000;
LUT4 lut_inst_1595 (
  .F(lut_f_1595),
  .I0(lut_f_1592),
  .I1(lut_f_1593),
  .I2(lut_f_1594),
  .I3(gw_vcc)
);
defparam lut_inst_1595.INIT = 16'h8000;
LUT4 lut_inst_1596 (
  .F(lut_f_1596),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1596.INIT = 16'h8000;
LUT4 lut_inst_1597 (
  .F(lut_f_1597),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1597.INIT = 16'h8000;
LUT4 lut_inst_1598 (
  .F(lut_f_1598),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1598.INIT = 16'h8000;
LUT4 lut_inst_1599 (
  .F(lut_f_1599),
  .I0(lut_f_1596),
  .I1(lut_f_1597),
  .I2(lut_f_1598),
  .I3(gw_vcc)
);
defparam lut_inst_1599.INIT = 16'h8000;
LUT4 lut_inst_1600 (
  .F(lut_f_1600),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1600.INIT = 16'h8000;
LUT4 lut_inst_1601 (
  .F(lut_f_1601),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1601.INIT = 16'h8000;
LUT4 lut_inst_1602 (
  .F(lut_f_1602),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1602.INIT = 16'h8000;
LUT4 lut_inst_1603 (
  .F(lut_f_1603),
  .I0(lut_f_1600),
  .I1(lut_f_1601),
  .I2(lut_f_1602),
  .I3(gw_vcc)
);
defparam lut_inst_1603.INIT = 16'h8000;
LUT4 lut_inst_1604 (
  .F(lut_f_1604),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1604.INIT = 16'h8000;
LUT4 lut_inst_1605 (
  .F(lut_f_1605),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1605.INIT = 16'h8000;
LUT4 lut_inst_1606 (
  .F(lut_f_1606),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1606.INIT = 16'h8000;
LUT4 lut_inst_1607 (
  .F(lut_f_1607),
  .I0(lut_f_1604),
  .I1(lut_f_1605),
  .I2(lut_f_1606),
  .I3(gw_vcc)
);
defparam lut_inst_1607.INIT = 16'h8000;
LUT4 lut_inst_1608 (
  .F(lut_f_1608),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1608.INIT = 16'h8000;
LUT4 lut_inst_1609 (
  .F(lut_f_1609),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1609.INIT = 16'h8000;
LUT4 lut_inst_1610 (
  .F(lut_f_1610),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1610.INIT = 16'h8000;
LUT4 lut_inst_1611 (
  .F(lut_f_1611),
  .I0(lut_f_1608),
  .I1(lut_f_1609),
  .I2(lut_f_1610),
  .I3(gw_vcc)
);
defparam lut_inst_1611.INIT = 16'h8000;
LUT4 lut_inst_1612 (
  .F(lut_f_1612),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1612.INIT = 16'h8000;
LUT4 lut_inst_1613 (
  .F(lut_f_1613),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1613.INIT = 16'h8000;
LUT4 lut_inst_1614 (
  .F(lut_f_1614),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1614.INIT = 16'h8000;
LUT4 lut_inst_1615 (
  .F(lut_f_1615),
  .I0(lut_f_1612),
  .I1(lut_f_1613),
  .I2(lut_f_1614),
  .I3(gw_vcc)
);
defparam lut_inst_1615.INIT = 16'h8000;
LUT4 lut_inst_1616 (
  .F(lut_f_1616),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1616.INIT = 16'h8000;
LUT4 lut_inst_1617 (
  .F(lut_f_1617),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1617.INIT = 16'h8000;
LUT4 lut_inst_1618 (
  .F(lut_f_1618),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1618.INIT = 16'h8000;
LUT4 lut_inst_1619 (
  .F(lut_f_1619),
  .I0(lut_f_1616),
  .I1(lut_f_1617),
  .I2(lut_f_1618),
  .I3(gw_vcc)
);
defparam lut_inst_1619.INIT = 16'h8000;
LUT4 lut_inst_1620 (
  .F(lut_f_1620),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1620.INIT = 16'h8000;
LUT4 lut_inst_1621 (
  .F(lut_f_1621),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1621.INIT = 16'h8000;
LUT4 lut_inst_1622 (
  .F(lut_f_1622),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1622.INIT = 16'h8000;
LUT4 lut_inst_1623 (
  .F(lut_f_1623),
  .I0(lut_f_1620),
  .I1(lut_f_1621),
  .I2(lut_f_1622),
  .I3(gw_vcc)
);
defparam lut_inst_1623.INIT = 16'h8000;
LUT4 lut_inst_1624 (
  .F(lut_f_1624),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1624.INIT = 16'h8000;
LUT4 lut_inst_1625 (
  .F(lut_f_1625),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1625.INIT = 16'h8000;
LUT4 lut_inst_1626 (
  .F(lut_f_1626),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1626.INIT = 16'h8000;
LUT4 lut_inst_1627 (
  .F(lut_f_1627),
  .I0(lut_f_1624),
  .I1(lut_f_1625),
  .I2(lut_f_1626),
  .I3(gw_vcc)
);
defparam lut_inst_1627.INIT = 16'h8000;
LUT4 lut_inst_1628 (
  .F(lut_f_1628),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1628.INIT = 16'h8000;
LUT4 lut_inst_1629 (
  .F(lut_f_1629),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1629.INIT = 16'h8000;
LUT4 lut_inst_1630 (
  .F(lut_f_1630),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1630.INIT = 16'h8000;
LUT4 lut_inst_1631 (
  .F(lut_f_1631),
  .I0(lut_f_1628),
  .I1(lut_f_1629),
  .I2(lut_f_1630),
  .I3(gw_vcc)
);
defparam lut_inst_1631.INIT = 16'h8000;
LUT4 lut_inst_1632 (
  .F(lut_f_1632),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1632.INIT = 16'h8000;
LUT4 lut_inst_1633 (
  .F(lut_f_1633),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1633.INIT = 16'h8000;
LUT4 lut_inst_1634 (
  .F(lut_f_1634),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1634.INIT = 16'h8000;
LUT4 lut_inst_1635 (
  .F(lut_f_1635),
  .I0(lut_f_1632),
  .I1(lut_f_1633),
  .I2(lut_f_1634),
  .I3(gw_vcc)
);
defparam lut_inst_1635.INIT = 16'h8000;
LUT4 lut_inst_1636 (
  .F(lut_f_1636),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1636.INIT = 16'h8000;
LUT4 lut_inst_1637 (
  .F(lut_f_1637),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1637.INIT = 16'h8000;
LUT4 lut_inst_1638 (
  .F(lut_f_1638),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1638.INIT = 16'h8000;
LUT4 lut_inst_1639 (
  .F(lut_f_1639),
  .I0(lut_f_1636),
  .I1(lut_f_1637),
  .I2(lut_f_1638),
  .I3(gw_vcc)
);
defparam lut_inst_1639.INIT = 16'h8000;
LUT4 lut_inst_1640 (
  .F(lut_f_1640),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1640.INIT = 16'h8000;
LUT4 lut_inst_1641 (
  .F(lut_f_1641),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1641.INIT = 16'h8000;
LUT4 lut_inst_1642 (
  .F(lut_f_1642),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1642.INIT = 16'h8000;
LUT4 lut_inst_1643 (
  .F(lut_f_1643),
  .I0(lut_f_1640),
  .I1(lut_f_1641),
  .I2(lut_f_1642),
  .I3(gw_vcc)
);
defparam lut_inst_1643.INIT = 16'h8000;
LUT4 lut_inst_1644 (
  .F(lut_f_1644),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1644.INIT = 16'h8000;
LUT4 lut_inst_1645 (
  .F(lut_f_1645),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1645.INIT = 16'h8000;
LUT4 lut_inst_1646 (
  .F(lut_f_1646),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1646.INIT = 16'h8000;
LUT4 lut_inst_1647 (
  .F(lut_f_1647),
  .I0(lut_f_1644),
  .I1(lut_f_1645),
  .I2(lut_f_1646),
  .I3(gw_vcc)
);
defparam lut_inst_1647.INIT = 16'h8000;
LUT4 lut_inst_1648 (
  .F(lut_f_1648),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1648.INIT = 16'h8000;
LUT4 lut_inst_1649 (
  .F(lut_f_1649),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1649.INIT = 16'h8000;
LUT4 lut_inst_1650 (
  .F(lut_f_1650),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1650.INIT = 16'h8000;
LUT4 lut_inst_1651 (
  .F(lut_f_1651),
  .I0(lut_f_1648),
  .I1(lut_f_1649),
  .I2(lut_f_1650),
  .I3(gw_vcc)
);
defparam lut_inst_1651.INIT = 16'h8000;
LUT4 lut_inst_1652 (
  .F(lut_f_1652),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1652.INIT = 16'h8000;
LUT4 lut_inst_1653 (
  .F(lut_f_1653),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1653.INIT = 16'h8000;
LUT4 lut_inst_1654 (
  .F(lut_f_1654),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1654.INIT = 16'h8000;
LUT4 lut_inst_1655 (
  .F(lut_f_1655),
  .I0(lut_f_1652),
  .I1(lut_f_1653),
  .I2(lut_f_1654),
  .I3(gw_vcc)
);
defparam lut_inst_1655.INIT = 16'h8000;
LUT4 lut_inst_1656 (
  .F(lut_f_1656),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1656.INIT = 16'h8000;
LUT4 lut_inst_1657 (
  .F(lut_f_1657),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1657.INIT = 16'h8000;
LUT4 lut_inst_1658 (
  .F(lut_f_1658),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1658.INIT = 16'h8000;
LUT4 lut_inst_1659 (
  .F(lut_f_1659),
  .I0(lut_f_1656),
  .I1(lut_f_1657),
  .I2(lut_f_1658),
  .I3(gw_vcc)
);
defparam lut_inst_1659.INIT = 16'h8000;
LUT4 lut_inst_1660 (
  .F(lut_f_1660),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1660.INIT = 16'h8000;
LUT4 lut_inst_1661 (
  .F(lut_f_1661),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_1661.INIT = 16'h8000;
LUT4 lut_inst_1662 (
  .F(lut_f_1662),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1662.INIT = 16'h8000;
LUT4 lut_inst_1663 (
  .F(lut_f_1663),
  .I0(lut_f_1660),
  .I1(lut_f_1661),
  .I2(lut_f_1662),
  .I3(gw_vcc)
);
defparam lut_inst_1663.INIT = 16'h8000;
LUT4 lut_inst_1664 (
  .F(lut_f_1664),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1664.INIT = 16'h8000;
LUT4 lut_inst_1665 (
  .F(lut_f_1665),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1665.INIT = 16'h8000;
LUT4 lut_inst_1666 (
  .F(lut_f_1666),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1666.INIT = 16'h8000;
LUT4 lut_inst_1667 (
  .F(lut_f_1667),
  .I0(lut_f_1664),
  .I1(lut_f_1665),
  .I2(lut_f_1666),
  .I3(gw_vcc)
);
defparam lut_inst_1667.INIT = 16'h8000;
LUT4 lut_inst_1668 (
  .F(lut_f_1668),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1668.INIT = 16'h8000;
LUT4 lut_inst_1669 (
  .F(lut_f_1669),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1669.INIT = 16'h8000;
LUT4 lut_inst_1670 (
  .F(lut_f_1670),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1670.INIT = 16'h8000;
LUT4 lut_inst_1671 (
  .F(lut_f_1671),
  .I0(lut_f_1668),
  .I1(lut_f_1669),
  .I2(lut_f_1670),
  .I3(gw_vcc)
);
defparam lut_inst_1671.INIT = 16'h8000;
LUT4 lut_inst_1672 (
  .F(lut_f_1672),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1672.INIT = 16'h8000;
LUT4 lut_inst_1673 (
  .F(lut_f_1673),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1673.INIT = 16'h8000;
LUT4 lut_inst_1674 (
  .F(lut_f_1674),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1674.INIT = 16'h8000;
LUT4 lut_inst_1675 (
  .F(lut_f_1675),
  .I0(lut_f_1672),
  .I1(lut_f_1673),
  .I2(lut_f_1674),
  .I3(gw_vcc)
);
defparam lut_inst_1675.INIT = 16'h8000;
LUT4 lut_inst_1676 (
  .F(lut_f_1676),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1676.INIT = 16'h8000;
LUT4 lut_inst_1677 (
  .F(lut_f_1677),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1677.INIT = 16'h8000;
LUT4 lut_inst_1678 (
  .F(lut_f_1678),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1678.INIT = 16'h8000;
LUT4 lut_inst_1679 (
  .F(lut_f_1679),
  .I0(lut_f_1676),
  .I1(lut_f_1677),
  .I2(lut_f_1678),
  .I3(gw_vcc)
);
defparam lut_inst_1679.INIT = 16'h8000;
LUT4 lut_inst_1680 (
  .F(lut_f_1680),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1680.INIT = 16'h8000;
LUT4 lut_inst_1681 (
  .F(lut_f_1681),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1681.INIT = 16'h8000;
LUT4 lut_inst_1682 (
  .F(lut_f_1682),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1682.INIT = 16'h8000;
LUT4 lut_inst_1683 (
  .F(lut_f_1683),
  .I0(lut_f_1680),
  .I1(lut_f_1681),
  .I2(lut_f_1682),
  .I3(gw_vcc)
);
defparam lut_inst_1683.INIT = 16'h8000;
LUT4 lut_inst_1684 (
  .F(lut_f_1684),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1684.INIT = 16'h8000;
LUT4 lut_inst_1685 (
  .F(lut_f_1685),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1685.INIT = 16'h8000;
LUT4 lut_inst_1686 (
  .F(lut_f_1686),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1686.INIT = 16'h8000;
LUT4 lut_inst_1687 (
  .F(lut_f_1687),
  .I0(lut_f_1684),
  .I1(lut_f_1685),
  .I2(lut_f_1686),
  .I3(gw_vcc)
);
defparam lut_inst_1687.INIT = 16'h8000;
LUT4 lut_inst_1688 (
  .F(lut_f_1688),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1688.INIT = 16'h8000;
LUT4 lut_inst_1689 (
  .F(lut_f_1689),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1689.INIT = 16'h8000;
LUT4 lut_inst_1690 (
  .F(lut_f_1690),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1690.INIT = 16'h8000;
LUT4 lut_inst_1691 (
  .F(lut_f_1691),
  .I0(lut_f_1688),
  .I1(lut_f_1689),
  .I2(lut_f_1690),
  .I3(gw_vcc)
);
defparam lut_inst_1691.INIT = 16'h8000;
LUT4 lut_inst_1692 (
  .F(lut_f_1692),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1692.INIT = 16'h8000;
LUT4 lut_inst_1693 (
  .F(lut_f_1693),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1693.INIT = 16'h8000;
LUT4 lut_inst_1694 (
  .F(lut_f_1694),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1694.INIT = 16'h8000;
LUT4 lut_inst_1695 (
  .F(lut_f_1695),
  .I0(lut_f_1692),
  .I1(lut_f_1693),
  .I2(lut_f_1694),
  .I3(gw_vcc)
);
defparam lut_inst_1695.INIT = 16'h8000;
LUT4 lut_inst_1696 (
  .F(lut_f_1696),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1696.INIT = 16'h8000;
LUT4 lut_inst_1697 (
  .F(lut_f_1697),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1697.INIT = 16'h8000;
LUT4 lut_inst_1698 (
  .F(lut_f_1698),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1698.INIT = 16'h8000;
LUT4 lut_inst_1699 (
  .F(lut_f_1699),
  .I0(lut_f_1696),
  .I1(lut_f_1697),
  .I2(lut_f_1698),
  .I3(gw_vcc)
);
defparam lut_inst_1699.INIT = 16'h8000;
LUT4 lut_inst_1700 (
  .F(lut_f_1700),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1700.INIT = 16'h8000;
LUT4 lut_inst_1701 (
  .F(lut_f_1701),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1701.INIT = 16'h8000;
LUT4 lut_inst_1702 (
  .F(lut_f_1702),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1702.INIT = 16'h8000;
LUT4 lut_inst_1703 (
  .F(lut_f_1703),
  .I0(lut_f_1700),
  .I1(lut_f_1701),
  .I2(lut_f_1702),
  .I3(gw_vcc)
);
defparam lut_inst_1703.INIT = 16'h8000;
LUT4 lut_inst_1704 (
  .F(lut_f_1704),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1704.INIT = 16'h8000;
LUT4 lut_inst_1705 (
  .F(lut_f_1705),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1705.INIT = 16'h8000;
LUT4 lut_inst_1706 (
  .F(lut_f_1706),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1706.INIT = 16'h8000;
LUT4 lut_inst_1707 (
  .F(lut_f_1707),
  .I0(lut_f_1704),
  .I1(lut_f_1705),
  .I2(lut_f_1706),
  .I3(gw_vcc)
);
defparam lut_inst_1707.INIT = 16'h8000;
LUT4 lut_inst_1708 (
  .F(lut_f_1708),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1708.INIT = 16'h8000;
LUT4 lut_inst_1709 (
  .F(lut_f_1709),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1709.INIT = 16'h8000;
LUT4 lut_inst_1710 (
  .F(lut_f_1710),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1710.INIT = 16'h8000;
LUT4 lut_inst_1711 (
  .F(lut_f_1711),
  .I0(lut_f_1708),
  .I1(lut_f_1709),
  .I2(lut_f_1710),
  .I3(gw_vcc)
);
defparam lut_inst_1711.INIT = 16'h8000;
LUT4 lut_inst_1712 (
  .F(lut_f_1712),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1712.INIT = 16'h8000;
LUT4 lut_inst_1713 (
  .F(lut_f_1713),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1713.INIT = 16'h8000;
LUT4 lut_inst_1714 (
  .F(lut_f_1714),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1714.INIT = 16'h8000;
LUT4 lut_inst_1715 (
  .F(lut_f_1715),
  .I0(lut_f_1712),
  .I1(lut_f_1713),
  .I2(lut_f_1714),
  .I3(gw_vcc)
);
defparam lut_inst_1715.INIT = 16'h8000;
LUT4 lut_inst_1716 (
  .F(lut_f_1716),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1716.INIT = 16'h8000;
LUT4 lut_inst_1717 (
  .F(lut_f_1717),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1717.INIT = 16'h8000;
LUT4 lut_inst_1718 (
  .F(lut_f_1718),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1718.INIT = 16'h8000;
LUT4 lut_inst_1719 (
  .F(lut_f_1719),
  .I0(lut_f_1716),
  .I1(lut_f_1717),
  .I2(lut_f_1718),
  .I3(gw_vcc)
);
defparam lut_inst_1719.INIT = 16'h8000;
LUT4 lut_inst_1720 (
  .F(lut_f_1720),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1720.INIT = 16'h8000;
LUT4 lut_inst_1721 (
  .F(lut_f_1721),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1721.INIT = 16'h8000;
LUT4 lut_inst_1722 (
  .F(lut_f_1722),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1722.INIT = 16'h8000;
LUT4 lut_inst_1723 (
  .F(lut_f_1723),
  .I0(lut_f_1720),
  .I1(lut_f_1721),
  .I2(lut_f_1722),
  .I3(gw_vcc)
);
defparam lut_inst_1723.INIT = 16'h8000;
LUT4 lut_inst_1724 (
  .F(lut_f_1724),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1724.INIT = 16'h8000;
LUT4 lut_inst_1725 (
  .F(lut_f_1725),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1725.INIT = 16'h8000;
LUT4 lut_inst_1726 (
  .F(lut_f_1726),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1726.INIT = 16'h8000;
LUT4 lut_inst_1727 (
  .F(lut_f_1727),
  .I0(lut_f_1724),
  .I1(lut_f_1725),
  .I2(lut_f_1726),
  .I3(gw_vcc)
);
defparam lut_inst_1727.INIT = 16'h8000;
LUT4 lut_inst_1728 (
  .F(lut_f_1728),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1728.INIT = 16'h8000;
LUT4 lut_inst_1729 (
  .F(lut_f_1729),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1729.INIT = 16'h8000;
LUT4 lut_inst_1730 (
  .F(lut_f_1730),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1730.INIT = 16'h8000;
LUT4 lut_inst_1731 (
  .F(lut_f_1731),
  .I0(lut_f_1728),
  .I1(lut_f_1729),
  .I2(lut_f_1730),
  .I3(gw_vcc)
);
defparam lut_inst_1731.INIT = 16'h8000;
LUT4 lut_inst_1732 (
  .F(lut_f_1732),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1732.INIT = 16'h8000;
LUT4 lut_inst_1733 (
  .F(lut_f_1733),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1733.INIT = 16'h8000;
LUT4 lut_inst_1734 (
  .F(lut_f_1734),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1734.INIT = 16'h8000;
LUT4 lut_inst_1735 (
  .F(lut_f_1735),
  .I0(lut_f_1732),
  .I1(lut_f_1733),
  .I2(lut_f_1734),
  .I3(gw_vcc)
);
defparam lut_inst_1735.INIT = 16'h8000;
LUT4 lut_inst_1736 (
  .F(lut_f_1736),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1736.INIT = 16'h8000;
LUT4 lut_inst_1737 (
  .F(lut_f_1737),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1737.INIT = 16'h8000;
LUT4 lut_inst_1738 (
  .F(lut_f_1738),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1738.INIT = 16'h8000;
LUT4 lut_inst_1739 (
  .F(lut_f_1739),
  .I0(lut_f_1736),
  .I1(lut_f_1737),
  .I2(lut_f_1738),
  .I3(gw_vcc)
);
defparam lut_inst_1739.INIT = 16'h8000;
LUT4 lut_inst_1740 (
  .F(lut_f_1740),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1740.INIT = 16'h8000;
LUT4 lut_inst_1741 (
  .F(lut_f_1741),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1741.INIT = 16'h8000;
LUT4 lut_inst_1742 (
  .F(lut_f_1742),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1742.INIT = 16'h8000;
LUT4 lut_inst_1743 (
  .F(lut_f_1743),
  .I0(lut_f_1740),
  .I1(lut_f_1741),
  .I2(lut_f_1742),
  .I3(gw_vcc)
);
defparam lut_inst_1743.INIT = 16'h8000;
LUT4 lut_inst_1744 (
  .F(lut_f_1744),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1744.INIT = 16'h8000;
LUT4 lut_inst_1745 (
  .F(lut_f_1745),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1745.INIT = 16'h8000;
LUT4 lut_inst_1746 (
  .F(lut_f_1746),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1746.INIT = 16'h8000;
LUT4 lut_inst_1747 (
  .F(lut_f_1747),
  .I0(lut_f_1744),
  .I1(lut_f_1745),
  .I2(lut_f_1746),
  .I3(gw_vcc)
);
defparam lut_inst_1747.INIT = 16'h8000;
LUT4 lut_inst_1748 (
  .F(lut_f_1748),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1748.INIT = 16'h8000;
LUT4 lut_inst_1749 (
  .F(lut_f_1749),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1749.INIT = 16'h8000;
LUT4 lut_inst_1750 (
  .F(lut_f_1750),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1750.INIT = 16'h8000;
LUT4 lut_inst_1751 (
  .F(lut_f_1751),
  .I0(lut_f_1748),
  .I1(lut_f_1749),
  .I2(lut_f_1750),
  .I3(gw_vcc)
);
defparam lut_inst_1751.INIT = 16'h8000;
LUT4 lut_inst_1752 (
  .F(lut_f_1752),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1752.INIT = 16'h8000;
LUT4 lut_inst_1753 (
  .F(lut_f_1753),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1753.INIT = 16'h8000;
LUT4 lut_inst_1754 (
  .F(lut_f_1754),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1754.INIT = 16'h8000;
LUT4 lut_inst_1755 (
  .F(lut_f_1755),
  .I0(lut_f_1752),
  .I1(lut_f_1753),
  .I2(lut_f_1754),
  .I3(gw_vcc)
);
defparam lut_inst_1755.INIT = 16'h8000;
LUT4 lut_inst_1756 (
  .F(lut_f_1756),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1756.INIT = 16'h8000;
LUT4 lut_inst_1757 (
  .F(lut_f_1757),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1757.INIT = 16'h8000;
LUT4 lut_inst_1758 (
  .F(lut_f_1758),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1758.INIT = 16'h8000;
LUT4 lut_inst_1759 (
  .F(lut_f_1759),
  .I0(lut_f_1756),
  .I1(lut_f_1757),
  .I2(lut_f_1758),
  .I3(gw_vcc)
);
defparam lut_inst_1759.INIT = 16'h8000;
LUT4 lut_inst_1760 (
  .F(lut_f_1760),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1760.INIT = 16'h8000;
LUT4 lut_inst_1761 (
  .F(lut_f_1761),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1761.INIT = 16'h8000;
LUT4 lut_inst_1762 (
  .F(lut_f_1762),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1762.INIT = 16'h8000;
LUT4 lut_inst_1763 (
  .F(lut_f_1763),
  .I0(lut_f_1760),
  .I1(lut_f_1761),
  .I2(lut_f_1762),
  .I3(gw_vcc)
);
defparam lut_inst_1763.INIT = 16'h8000;
LUT4 lut_inst_1764 (
  .F(lut_f_1764),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1764.INIT = 16'h8000;
LUT4 lut_inst_1765 (
  .F(lut_f_1765),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1765.INIT = 16'h8000;
LUT4 lut_inst_1766 (
  .F(lut_f_1766),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1766.INIT = 16'h8000;
LUT4 lut_inst_1767 (
  .F(lut_f_1767),
  .I0(lut_f_1764),
  .I1(lut_f_1765),
  .I2(lut_f_1766),
  .I3(gw_vcc)
);
defparam lut_inst_1767.INIT = 16'h8000;
LUT4 lut_inst_1768 (
  .F(lut_f_1768),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1768.INIT = 16'h8000;
LUT4 lut_inst_1769 (
  .F(lut_f_1769),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1769.INIT = 16'h8000;
LUT4 lut_inst_1770 (
  .F(lut_f_1770),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1770.INIT = 16'h8000;
LUT4 lut_inst_1771 (
  .F(lut_f_1771),
  .I0(lut_f_1768),
  .I1(lut_f_1769),
  .I2(lut_f_1770),
  .I3(gw_vcc)
);
defparam lut_inst_1771.INIT = 16'h8000;
LUT4 lut_inst_1772 (
  .F(lut_f_1772),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1772.INIT = 16'h8000;
LUT4 lut_inst_1773 (
  .F(lut_f_1773),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1773.INIT = 16'h8000;
LUT4 lut_inst_1774 (
  .F(lut_f_1774),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1774.INIT = 16'h8000;
LUT4 lut_inst_1775 (
  .F(lut_f_1775),
  .I0(lut_f_1772),
  .I1(lut_f_1773),
  .I2(lut_f_1774),
  .I3(gw_vcc)
);
defparam lut_inst_1775.INIT = 16'h8000;
LUT4 lut_inst_1776 (
  .F(lut_f_1776),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1776.INIT = 16'h8000;
LUT4 lut_inst_1777 (
  .F(lut_f_1777),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1777.INIT = 16'h8000;
LUT4 lut_inst_1778 (
  .F(lut_f_1778),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1778.INIT = 16'h8000;
LUT4 lut_inst_1779 (
  .F(lut_f_1779),
  .I0(lut_f_1776),
  .I1(lut_f_1777),
  .I2(lut_f_1778),
  .I3(gw_vcc)
);
defparam lut_inst_1779.INIT = 16'h8000;
LUT4 lut_inst_1780 (
  .F(lut_f_1780),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1780.INIT = 16'h8000;
LUT4 lut_inst_1781 (
  .F(lut_f_1781),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1781.INIT = 16'h8000;
LUT4 lut_inst_1782 (
  .F(lut_f_1782),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1782.INIT = 16'h8000;
LUT4 lut_inst_1783 (
  .F(lut_f_1783),
  .I0(lut_f_1780),
  .I1(lut_f_1781),
  .I2(lut_f_1782),
  .I3(gw_vcc)
);
defparam lut_inst_1783.INIT = 16'h8000;
LUT4 lut_inst_1784 (
  .F(lut_f_1784),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1784.INIT = 16'h8000;
LUT4 lut_inst_1785 (
  .F(lut_f_1785),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1785.INIT = 16'h8000;
LUT4 lut_inst_1786 (
  .F(lut_f_1786),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1786.INIT = 16'h8000;
LUT4 lut_inst_1787 (
  .F(lut_f_1787),
  .I0(lut_f_1784),
  .I1(lut_f_1785),
  .I2(lut_f_1786),
  .I3(gw_vcc)
);
defparam lut_inst_1787.INIT = 16'h8000;
LUT4 lut_inst_1788 (
  .F(lut_f_1788),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1788.INIT = 16'h8000;
LUT4 lut_inst_1789 (
  .F(lut_f_1789),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_1789.INIT = 16'h8000;
LUT4 lut_inst_1790 (
  .F(lut_f_1790),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1790.INIT = 16'h8000;
LUT4 lut_inst_1791 (
  .F(lut_f_1791),
  .I0(lut_f_1788),
  .I1(lut_f_1789),
  .I2(lut_f_1790),
  .I3(gw_vcc)
);
defparam lut_inst_1791.INIT = 16'h8000;
LUT4 lut_inst_1792 (
  .F(lut_f_1792),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1792.INIT = 16'h8000;
LUT4 lut_inst_1793 (
  .F(lut_f_1793),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1793.INIT = 16'h8000;
LUT4 lut_inst_1794 (
  .F(lut_f_1794),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1794.INIT = 16'h8000;
LUT4 lut_inst_1795 (
  .F(lut_f_1795),
  .I0(lut_f_1792),
  .I1(lut_f_1793),
  .I2(lut_f_1794),
  .I3(gw_vcc)
);
defparam lut_inst_1795.INIT = 16'h8000;
LUT4 lut_inst_1796 (
  .F(lut_f_1796),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1796.INIT = 16'h8000;
LUT4 lut_inst_1797 (
  .F(lut_f_1797),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1797.INIT = 16'h8000;
LUT4 lut_inst_1798 (
  .F(lut_f_1798),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1798.INIT = 16'h8000;
LUT4 lut_inst_1799 (
  .F(lut_f_1799),
  .I0(lut_f_1796),
  .I1(lut_f_1797),
  .I2(lut_f_1798),
  .I3(gw_vcc)
);
defparam lut_inst_1799.INIT = 16'h8000;
LUT4 lut_inst_1800 (
  .F(lut_f_1800),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1800.INIT = 16'h8000;
LUT4 lut_inst_1801 (
  .F(lut_f_1801),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1801.INIT = 16'h8000;
LUT4 lut_inst_1802 (
  .F(lut_f_1802),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1802.INIT = 16'h8000;
LUT4 lut_inst_1803 (
  .F(lut_f_1803),
  .I0(lut_f_1800),
  .I1(lut_f_1801),
  .I2(lut_f_1802),
  .I3(gw_vcc)
);
defparam lut_inst_1803.INIT = 16'h8000;
LUT4 lut_inst_1804 (
  .F(lut_f_1804),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1804.INIT = 16'h8000;
LUT4 lut_inst_1805 (
  .F(lut_f_1805),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1805.INIT = 16'h8000;
LUT4 lut_inst_1806 (
  .F(lut_f_1806),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1806.INIT = 16'h8000;
LUT4 lut_inst_1807 (
  .F(lut_f_1807),
  .I0(lut_f_1804),
  .I1(lut_f_1805),
  .I2(lut_f_1806),
  .I3(gw_vcc)
);
defparam lut_inst_1807.INIT = 16'h8000;
LUT4 lut_inst_1808 (
  .F(lut_f_1808),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1808.INIT = 16'h8000;
LUT4 lut_inst_1809 (
  .F(lut_f_1809),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1809.INIT = 16'h8000;
LUT4 lut_inst_1810 (
  .F(lut_f_1810),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1810.INIT = 16'h8000;
LUT4 lut_inst_1811 (
  .F(lut_f_1811),
  .I0(lut_f_1808),
  .I1(lut_f_1809),
  .I2(lut_f_1810),
  .I3(gw_vcc)
);
defparam lut_inst_1811.INIT = 16'h8000;
LUT4 lut_inst_1812 (
  .F(lut_f_1812),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1812.INIT = 16'h8000;
LUT4 lut_inst_1813 (
  .F(lut_f_1813),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1813.INIT = 16'h8000;
LUT4 lut_inst_1814 (
  .F(lut_f_1814),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1814.INIT = 16'h8000;
LUT4 lut_inst_1815 (
  .F(lut_f_1815),
  .I0(lut_f_1812),
  .I1(lut_f_1813),
  .I2(lut_f_1814),
  .I3(gw_vcc)
);
defparam lut_inst_1815.INIT = 16'h8000;
LUT4 lut_inst_1816 (
  .F(lut_f_1816),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1816.INIT = 16'h8000;
LUT4 lut_inst_1817 (
  .F(lut_f_1817),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1817.INIT = 16'h8000;
LUT4 lut_inst_1818 (
  .F(lut_f_1818),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1818.INIT = 16'h8000;
LUT4 lut_inst_1819 (
  .F(lut_f_1819),
  .I0(lut_f_1816),
  .I1(lut_f_1817),
  .I2(lut_f_1818),
  .I3(gw_vcc)
);
defparam lut_inst_1819.INIT = 16'h8000;
LUT4 lut_inst_1820 (
  .F(lut_f_1820),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1820.INIT = 16'h8000;
LUT4 lut_inst_1821 (
  .F(lut_f_1821),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1821.INIT = 16'h8000;
LUT4 lut_inst_1822 (
  .F(lut_f_1822),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1822.INIT = 16'h8000;
LUT4 lut_inst_1823 (
  .F(lut_f_1823),
  .I0(lut_f_1820),
  .I1(lut_f_1821),
  .I2(lut_f_1822),
  .I3(gw_vcc)
);
defparam lut_inst_1823.INIT = 16'h8000;
LUT4 lut_inst_1824 (
  .F(lut_f_1824),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1824.INIT = 16'h8000;
LUT4 lut_inst_1825 (
  .F(lut_f_1825),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1825.INIT = 16'h8000;
LUT4 lut_inst_1826 (
  .F(lut_f_1826),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1826.INIT = 16'h8000;
LUT4 lut_inst_1827 (
  .F(lut_f_1827),
  .I0(lut_f_1824),
  .I1(lut_f_1825),
  .I2(lut_f_1826),
  .I3(gw_vcc)
);
defparam lut_inst_1827.INIT = 16'h8000;
LUT4 lut_inst_1828 (
  .F(lut_f_1828),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1828.INIT = 16'h8000;
LUT4 lut_inst_1829 (
  .F(lut_f_1829),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1829.INIT = 16'h8000;
LUT4 lut_inst_1830 (
  .F(lut_f_1830),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1830.INIT = 16'h8000;
LUT4 lut_inst_1831 (
  .F(lut_f_1831),
  .I0(lut_f_1828),
  .I1(lut_f_1829),
  .I2(lut_f_1830),
  .I3(gw_vcc)
);
defparam lut_inst_1831.INIT = 16'h8000;
LUT4 lut_inst_1832 (
  .F(lut_f_1832),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1832.INIT = 16'h8000;
LUT4 lut_inst_1833 (
  .F(lut_f_1833),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1833.INIT = 16'h8000;
LUT4 lut_inst_1834 (
  .F(lut_f_1834),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1834.INIT = 16'h8000;
LUT4 lut_inst_1835 (
  .F(lut_f_1835),
  .I0(lut_f_1832),
  .I1(lut_f_1833),
  .I2(lut_f_1834),
  .I3(gw_vcc)
);
defparam lut_inst_1835.INIT = 16'h8000;
LUT4 lut_inst_1836 (
  .F(lut_f_1836),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1836.INIT = 16'h8000;
LUT4 lut_inst_1837 (
  .F(lut_f_1837),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1837.INIT = 16'h8000;
LUT4 lut_inst_1838 (
  .F(lut_f_1838),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1838.INIT = 16'h8000;
LUT4 lut_inst_1839 (
  .F(lut_f_1839),
  .I0(lut_f_1836),
  .I1(lut_f_1837),
  .I2(lut_f_1838),
  .I3(gw_vcc)
);
defparam lut_inst_1839.INIT = 16'h8000;
LUT4 lut_inst_1840 (
  .F(lut_f_1840),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1840.INIT = 16'h8000;
LUT4 lut_inst_1841 (
  .F(lut_f_1841),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1841.INIT = 16'h8000;
LUT4 lut_inst_1842 (
  .F(lut_f_1842),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1842.INIT = 16'h8000;
LUT4 lut_inst_1843 (
  .F(lut_f_1843),
  .I0(lut_f_1840),
  .I1(lut_f_1841),
  .I2(lut_f_1842),
  .I3(gw_vcc)
);
defparam lut_inst_1843.INIT = 16'h8000;
LUT4 lut_inst_1844 (
  .F(lut_f_1844),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1844.INIT = 16'h8000;
LUT4 lut_inst_1845 (
  .F(lut_f_1845),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1845.INIT = 16'h8000;
LUT4 lut_inst_1846 (
  .F(lut_f_1846),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1846.INIT = 16'h8000;
LUT4 lut_inst_1847 (
  .F(lut_f_1847),
  .I0(lut_f_1844),
  .I1(lut_f_1845),
  .I2(lut_f_1846),
  .I3(gw_vcc)
);
defparam lut_inst_1847.INIT = 16'h8000;
LUT4 lut_inst_1848 (
  .F(lut_f_1848),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1848.INIT = 16'h8000;
LUT4 lut_inst_1849 (
  .F(lut_f_1849),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1849.INIT = 16'h8000;
LUT4 lut_inst_1850 (
  .F(lut_f_1850),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1850.INIT = 16'h8000;
LUT4 lut_inst_1851 (
  .F(lut_f_1851),
  .I0(lut_f_1848),
  .I1(lut_f_1849),
  .I2(lut_f_1850),
  .I3(gw_vcc)
);
defparam lut_inst_1851.INIT = 16'h8000;
LUT4 lut_inst_1852 (
  .F(lut_f_1852),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1852.INIT = 16'h8000;
LUT4 lut_inst_1853 (
  .F(lut_f_1853),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1853.INIT = 16'h8000;
LUT4 lut_inst_1854 (
  .F(lut_f_1854),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1854.INIT = 16'h8000;
LUT4 lut_inst_1855 (
  .F(lut_f_1855),
  .I0(lut_f_1852),
  .I1(lut_f_1853),
  .I2(lut_f_1854),
  .I3(gw_vcc)
);
defparam lut_inst_1855.INIT = 16'h8000;
LUT4 lut_inst_1856 (
  .F(lut_f_1856),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1856.INIT = 16'h8000;
LUT4 lut_inst_1857 (
  .F(lut_f_1857),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1857.INIT = 16'h8000;
LUT4 lut_inst_1858 (
  .F(lut_f_1858),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1858.INIT = 16'h8000;
LUT4 lut_inst_1859 (
  .F(lut_f_1859),
  .I0(lut_f_1856),
  .I1(lut_f_1857),
  .I2(lut_f_1858),
  .I3(gw_vcc)
);
defparam lut_inst_1859.INIT = 16'h8000;
LUT4 lut_inst_1860 (
  .F(lut_f_1860),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1860.INIT = 16'h8000;
LUT4 lut_inst_1861 (
  .F(lut_f_1861),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1861.INIT = 16'h8000;
LUT4 lut_inst_1862 (
  .F(lut_f_1862),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1862.INIT = 16'h8000;
LUT4 lut_inst_1863 (
  .F(lut_f_1863),
  .I0(lut_f_1860),
  .I1(lut_f_1861),
  .I2(lut_f_1862),
  .I3(gw_vcc)
);
defparam lut_inst_1863.INIT = 16'h8000;
LUT4 lut_inst_1864 (
  .F(lut_f_1864),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1864.INIT = 16'h8000;
LUT4 lut_inst_1865 (
  .F(lut_f_1865),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1865.INIT = 16'h8000;
LUT4 lut_inst_1866 (
  .F(lut_f_1866),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1866.INIT = 16'h8000;
LUT4 lut_inst_1867 (
  .F(lut_f_1867),
  .I0(lut_f_1864),
  .I1(lut_f_1865),
  .I2(lut_f_1866),
  .I3(gw_vcc)
);
defparam lut_inst_1867.INIT = 16'h8000;
LUT4 lut_inst_1868 (
  .F(lut_f_1868),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1868.INIT = 16'h8000;
LUT4 lut_inst_1869 (
  .F(lut_f_1869),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1869.INIT = 16'h8000;
LUT4 lut_inst_1870 (
  .F(lut_f_1870),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1870.INIT = 16'h8000;
LUT4 lut_inst_1871 (
  .F(lut_f_1871),
  .I0(lut_f_1868),
  .I1(lut_f_1869),
  .I2(lut_f_1870),
  .I3(gw_vcc)
);
defparam lut_inst_1871.INIT = 16'h8000;
LUT4 lut_inst_1872 (
  .F(lut_f_1872),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1872.INIT = 16'h8000;
LUT4 lut_inst_1873 (
  .F(lut_f_1873),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1873.INIT = 16'h8000;
LUT4 lut_inst_1874 (
  .F(lut_f_1874),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1874.INIT = 16'h8000;
LUT4 lut_inst_1875 (
  .F(lut_f_1875),
  .I0(lut_f_1872),
  .I1(lut_f_1873),
  .I2(lut_f_1874),
  .I3(gw_vcc)
);
defparam lut_inst_1875.INIT = 16'h8000;
LUT4 lut_inst_1876 (
  .F(lut_f_1876),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1876.INIT = 16'h8000;
LUT4 lut_inst_1877 (
  .F(lut_f_1877),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1877.INIT = 16'h8000;
LUT4 lut_inst_1878 (
  .F(lut_f_1878),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1878.INIT = 16'h8000;
LUT4 lut_inst_1879 (
  .F(lut_f_1879),
  .I0(lut_f_1876),
  .I1(lut_f_1877),
  .I2(lut_f_1878),
  .I3(gw_vcc)
);
defparam lut_inst_1879.INIT = 16'h8000;
LUT4 lut_inst_1880 (
  .F(lut_f_1880),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1880.INIT = 16'h8000;
LUT4 lut_inst_1881 (
  .F(lut_f_1881),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1881.INIT = 16'h8000;
LUT4 lut_inst_1882 (
  .F(lut_f_1882),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1882.INIT = 16'h8000;
LUT4 lut_inst_1883 (
  .F(lut_f_1883),
  .I0(lut_f_1880),
  .I1(lut_f_1881),
  .I2(lut_f_1882),
  .I3(gw_vcc)
);
defparam lut_inst_1883.INIT = 16'h8000;
LUT4 lut_inst_1884 (
  .F(lut_f_1884),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1884.INIT = 16'h8000;
LUT4 lut_inst_1885 (
  .F(lut_f_1885),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1885.INIT = 16'h8000;
LUT4 lut_inst_1886 (
  .F(lut_f_1886),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1886.INIT = 16'h8000;
LUT4 lut_inst_1887 (
  .F(lut_f_1887),
  .I0(lut_f_1884),
  .I1(lut_f_1885),
  .I2(lut_f_1886),
  .I3(gw_vcc)
);
defparam lut_inst_1887.INIT = 16'h8000;
LUT4 lut_inst_1888 (
  .F(lut_f_1888),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1888.INIT = 16'h8000;
LUT4 lut_inst_1889 (
  .F(lut_f_1889),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1889.INIT = 16'h8000;
LUT4 lut_inst_1890 (
  .F(lut_f_1890),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1890.INIT = 16'h8000;
LUT4 lut_inst_1891 (
  .F(lut_f_1891),
  .I0(lut_f_1888),
  .I1(lut_f_1889),
  .I2(lut_f_1890),
  .I3(gw_vcc)
);
defparam lut_inst_1891.INIT = 16'h8000;
LUT4 lut_inst_1892 (
  .F(lut_f_1892),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1892.INIT = 16'h8000;
LUT4 lut_inst_1893 (
  .F(lut_f_1893),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1893.INIT = 16'h8000;
LUT4 lut_inst_1894 (
  .F(lut_f_1894),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1894.INIT = 16'h8000;
LUT4 lut_inst_1895 (
  .F(lut_f_1895),
  .I0(lut_f_1892),
  .I1(lut_f_1893),
  .I2(lut_f_1894),
  .I3(gw_vcc)
);
defparam lut_inst_1895.INIT = 16'h8000;
LUT4 lut_inst_1896 (
  .F(lut_f_1896),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1896.INIT = 16'h8000;
LUT4 lut_inst_1897 (
  .F(lut_f_1897),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1897.INIT = 16'h8000;
LUT4 lut_inst_1898 (
  .F(lut_f_1898),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1898.INIT = 16'h8000;
LUT4 lut_inst_1899 (
  .F(lut_f_1899),
  .I0(lut_f_1896),
  .I1(lut_f_1897),
  .I2(lut_f_1898),
  .I3(gw_vcc)
);
defparam lut_inst_1899.INIT = 16'h8000;
LUT4 lut_inst_1900 (
  .F(lut_f_1900),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1900.INIT = 16'h8000;
LUT4 lut_inst_1901 (
  .F(lut_f_1901),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1901.INIT = 16'h8000;
LUT4 lut_inst_1902 (
  .F(lut_f_1902),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1902.INIT = 16'h8000;
LUT4 lut_inst_1903 (
  .F(lut_f_1903),
  .I0(lut_f_1900),
  .I1(lut_f_1901),
  .I2(lut_f_1902),
  .I3(gw_vcc)
);
defparam lut_inst_1903.INIT = 16'h8000;
LUT4 lut_inst_1904 (
  .F(lut_f_1904),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1904.INIT = 16'h8000;
LUT4 lut_inst_1905 (
  .F(lut_f_1905),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1905.INIT = 16'h8000;
LUT4 lut_inst_1906 (
  .F(lut_f_1906),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1906.INIT = 16'h8000;
LUT4 lut_inst_1907 (
  .F(lut_f_1907),
  .I0(lut_f_1904),
  .I1(lut_f_1905),
  .I2(lut_f_1906),
  .I3(gw_vcc)
);
defparam lut_inst_1907.INIT = 16'h8000;
LUT4 lut_inst_1908 (
  .F(lut_f_1908),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1908.INIT = 16'h8000;
LUT4 lut_inst_1909 (
  .F(lut_f_1909),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1909.INIT = 16'h8000;
LUT4 lut_inst_1910 (
  .F(lut_f_1910),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1910.INIT = 16'h8000;
LUT4 lut_inst_1911 (
  .F(lut_f_1911),
  .I0(lut_f_1908),
  .I1(lut_f_1909),
  .I2(lut_f_1910),
  .I3(gw_vcc)
);
defparam lut_inst_1911.INIT = 16'h8000;
LUT4 lut_inst_1912 (
  .F(lut_f_1912),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1912.INIT = 16'h8000;
LUT4 lut_inst_1913 (
  .F(lut_f_1913),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1913.INIT = 16'h8000;
LUT4 lut_inst_1914 (
  .F(lut_f_1914),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1914.INIT = 16'h8000;
LUT4 lut_inst_1915 (
  .F(lut_f_1915),
  .I0(lut_f_1912),
  .I1(lut_f_1913),
  .I2(lut_f_1914),
  .I3(gw_vcc)
);
defparam lut_inst_1915.INIT = 16'h8000;
LUT4 lut_inst_1916 (
  .F(lut_f_1916),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1916.INIT = 16'h8000;
LUT4 lut_inst_1917 (
  .F(lut_f_1917),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_1917.INIT = 16'h8000;
LUT4 lut_inst_1918 (
  .F(lut_f_1918),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1918.INIT = 16'h8000;
LUT4 lut_inst_1919 (
  .F(lut_f_1919),
  .I0(lut_f_1916),
  .I1(lut_f_1917),
  .I2(lut_f_1918),
  .I3(gw_vcc)
);
defparam lut_inst_1919.INIT = 16'h8000;
LUT4 lut_inst_1920 (
  .F(lut_f_1920),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1920.INIT = 16'h8000;
LUT4 lut_inst_1921 (
  .F(lut_f_1921),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1921.INIT = 16'h8000;
LUT4 lut_inst_1922 (
  .F(lut_f_1922),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1922.INIT = 16'h8000;
LUT4 lut_inst_1923 (
  .F(lut_f_1923),
  .I0(lut_f_1920),
  .I1(lut_f_1921),
  .I2(lut_f_1922),
  .I3(gw_vcc)
);
defparam lut_inst_1923.INIT = 16'h8000;
LUT4 lut_inst_1924 (
  .F(lut_f_1924),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1924.INIT = 16'h8000;
LUT4 lut_inst_1925 (
  .F(lut_f_1925),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1925.INIT = 16'h8000;
LUT4 lut_inst_1926 (
  .F(lut_f_1926),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1926.INIT = 16'h8000;
LUT4 lut_inst_1927 (
  .F(lut_f_1927),
  .I0(lut_f_1924),
  .I1(lut_f_1925),
  .I2(lut_f_1926),
  .I3(gw_vcc)
);
defparam lut_inst_1927.INIT = 16'h8000;
LUT4 lut_inst_1928 (
  .F(lut_f_1928),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1928.INIT = 16'h8000;
LUT4 lut_inst_1929 (
  .F(lut_f_1929),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1929.INIT = 16'h8000;
LUT4 lut_inst_1930 (
  .F(lut_f_1930),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1930.INIT = 16'h8000;
LUT4 lut_inst_1931 (
  .F(lut_f_1931),
  .I0(lut_f_1928),
  .I1(lut_f_1929),
  .I2(lut_f_1930),
  .I3(gw_vcc)
);
defparam lut_inst_1931.INIT = 16'h8000;
LUT4 lut_inst_1932 (
  .F(lut_f_1932),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1932.INIT = 16'h8000;
LUT4 lut_inst_1933 (
  .F(lut_f_1933),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1933.INIT = 16'h8000;
LUT4 lut_inst_1934 (
  .F(lut_f_1934),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1934.INIT = 16'h8000;
LUT4 lut_inst_1935 (
  .F(lut_f_1935),
  .I0(lut_f_1932),
  .I1(lut_f_1933),
  .I2(lut_f_1934),
  .I3(gw_vcc)
);
defparam lut_inst_1935.INIT = 16'h8000;
LUT4 lut_inst_1936 (
  .F(lut_f_1936),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1936.INIT = 16'h8000;
LUT4 lut_inst_1937 (
  .F(lut_f_1937),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1937.INIT = 16'h8000;
LUT4 lut_inst_1938 (
  .F(lut_f_1938),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1938.INIT = 16'h8000;
LUT4 lut_inst_1939 (
  .F(lut_f_1939),
  .I0(lut_f_1936),
  .I1(lut_f_1937),
  .I2(lut_f_1938),
  .I3(gw_vcc)
);
defparam lut_inst_1939.INIT = 16'h8000;
LUT4 lut_inst_1940 (
  .F(lut_f_1940),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1940.INIT = 16'h8000;
LUT4 lut_inst_1941 (
  .F(lut_f_1941),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1941.INIT = 16'h8000;
LUT4 lut_inst_1942 (
  .F(lut_f_1942),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1942.INIT = 16'h8000;
LUT4 lut_inst_1943 (
  .F(lut_f_1943),
  .I0(lut_f_1940),
  .I1(lut_f_1941),
  .I2(lut_f_1942),
  .I3(gw_vcc)
);
defparam lut_inst_1943.INIT = 16'h8000;
LUT4 lut_inst_1944 (
  .F(lut_f_1944),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1944.INIT = 16'h8000;
LUT4 lut_inst_1945 (
  .F(lut_f_1945),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1945.INIT = 16'h8000;
LUT4 lut_inst_1946 (
  .F(lut_f_1946),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1946.INIT = 16'h8000;
LUT4 lut_inst_1947 (
  .F(lut_f_1947),
  .I0(lut_f_1944),
  .I1(lut_f_1945),
  .I2(lut_f_1946),
  .I3(gw_vcc)
);
defparam lut_inst_1947.INIT = 16'h8000;
LUT4 lut_inst_1948 (
  .F(lut_f_1948),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1948.INIT = 16'h8000;
LUT4 lut_inst_1949 (
  .F(lut_f_1949),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1949.INIT = 16'h8000;
LUT4 lut_inst_1950 (
  .F(lut_f_1950),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1950.INIT = 16'h8000;
LUT4 lut_inst_1951 (
  .F(lut_f_1951),
  .I0(lut_f_1948),
  .I1(lut_f_1949),
  .I2(lut_f_1950),
  .I3(gw_vcc)
);
defparam lut_inst_1951.INIT = 16'h8000;
LUT4 lut_inst_1952 (
  .F(lut_f_1952),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1952.INIT = 16'h8000;
LUT4 lut_inst_1953 (
  .F(lut_f_1953),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1953.INIT = 16'h8000;
LUT4 lut_inst_1954 (
  .F(lut_f_1954),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1954.INIT = 16'h8000;
LUT4 lut_inst_1955 (
  .F(lut_f_1955),
  .I0(lut_f_1952),
  .I1(lut_f_1953),
  .I2(lut_f_1954),
  .I3(gw_vcc)
);
defparam lut_inst_1955.INIT = 16'h8000;
LUT4 lut_inst_1956 (
  .F(lut_f_1956),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1956.INIT = 16'h8000;
LUT4 lut_inst_1957 (
  .F(lut_f_1957),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1957.INIT = 16'h8000;
LUT4 lut_inst_1958 (
  .F(lut_f_1958),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1958.INIT = 16'h8000;
LUT4 lut_inst_1959 (
  .F(lut_f_1959),
  .I0(lut_f_1956),
  .I1(lut_f_1957),
  .I2(lut_f_1958),
  .I3(gw_vcc)
);
defparam lut_inst_1959.INIT = 16'h8000;
LUT4 lut_inst_1960 (
  .F(lut_f_1960),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1960.INIT = 16'h8000;
LUT4 lut_inst_1961 (
  .F(lut_f_1961),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1961.INIT = 16'h8000;
LUT4 lut_inst_1962 (
  .F(lut_f_1962),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1962.INIT = 16'h8000;
LUT4 lut_inst_1963 (
  .F(lut_f_1963),
  .I0(lut_f_1960),
  .I1(lut_f_1961),
  .I2(lut_f_1962),
  .I3(gw_vcc)
);
defparam lut_inst_1963.INIT = 16'h8000;
LUT4 lut_inst_1964 (
  .F(lut_f_1964),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1964.INIT = 16'h8000;
LUT4 lut_inst_1965 (
  .F(lut_f_1965),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1965.INIT = 16'h8000;
LUT4 lut_inst_1966 (
  .F(lut_f_1966),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1966.INIT = 16'h8000;
LUT4 lut_inst_1967 (
  .F(lut_f_1967),
  .I0(lut_f_1964),
  .I1(lut_f_1965),
  .I2(lut_f_1966),
  .I3(gw_vcc)
);
defparam lut_inst_1967.INIT = 16'h8000;
LUT4 lut_inst_1968 (
  .F(lut_f_1968),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1968.INIT = 16'h8000;
LUT4 lut_inst_1969 (
  .F(lut_f_1969),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1969.INIT = 16'h8000;
LUT4 lut_inst_1970 (
  .F(lut_f_1970),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1970.INIT = 16'h8000;
LUT4 lut_inst_1971 (
  .F(lut_f_1971),
  .I0(lut_f_1968),
  .I1(lut_f_1969),
  .I2(lut_f_1970),
  .I3(gw_vcc)
);
defparam lut_inst_1971.INIT = 16'h8000;
LUT4 lut_inst_1972 (
  .F(lut_f_1972),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_1972.INIT = 16'h8000;
LUT4 lut_inst_1973 (
  .F(lut_f_1973),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1973.INIT = 16'h8000;
LUT4 lut_inst_1974 (
  .F(lut_f_1974),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1974.INIT = 16'h8000;
LUT4 lut_inst_1975 (
  .F(lut_f_1975),
  .I0(lut_f_1972),
  .I1(lut_f_1973),
  .I2(lut_f_1974),
  .I3(gw_vcc)
);
defparam lut_inst_1975.INIT = 16'h8000;
LUT4 lut_inst_1976 (
  .F(lut_f_1976),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1976.INIT = 16'h8000;
LUT4 lut_inst_1977 (
  .F(lut_f_1977),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1977.INIT = 16'h8000;
LUT4 lut_inst_1978 (
  .F(lut_f_1978),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1978.INIT = 16'h8000;
LUT4 lut_inst_1979 (
  .F(lut_f_1979),
  .I0(lut_f_1976),
  .I1(lut_f_1977),
  .I2(lut_f_1978),
  .I3(gw_vcc)
);
defparam lut_inst_1979.INIT = 16'h8000;
LUT4 lut_inst_1980 (
  .F(lut_f_1980),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_1980.INIT = 16'h8000;
LUT4 lut_inst_1981 (
  .F(lut_f_1981),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1981.INIT = 16'h8000;
LUT4 lut_inst_1982 (
  .F(lut_f_1982),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1982.INIT = 16'h8000;
LUT4 lut_inst_1983 (
  .F(lut_f_1983),
  .I0(lut_f_1980),
  .I1(lut_f_1981),
  .I2(lut_f_1982),
  .I3(gw_vcc)
);
defparam lut_inst_1983.INIT = 16'h8000;
LUT4 lut_inst_1984 (
  .F(lut_f_1984),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1984.INIT = 16'h8000;
LUT4 lut_inst_1985 (
  .F(lut_f_1985),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1985.INIT = 16'h8000;
LUT4 lut_inst_1986 (
  .F(lut_f_1986),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1986.INIT = 16'h8000;
LUT4 lut_inst_1987 (
  .F(lut_f_1987),
  .I0(lut_f_1984),
  .I1(lut_f_1985),
  .I2(lut_f_1986),
  .I3(gw_vcc)
);
defparam lut_inst_1987.INIT = 16'h8000;
LUT4 lut_inst_1988 (
  .F(lut_f_1988),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_1988.INIT = 16'h8000;
LUT4 lut_inst_1989 (
  .F(lut_f_1989),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1989.INIT = 16'h8000;
LUT4 lut_inst_1990 (
  .F(lut_f_1990),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1990.INIT = 16'h8000;
LUT4 lut_inst_1991 (
  .F(lut_f_1991),
  .I0(lut_f_1988),
  .I1(lut_f_1989),
  .I2(lut_f_1990),
  .I3(gw_vcc)
);
defparam lut_inst_1991.INIT = 16'h8000;
LUT4 lut_inst_1992 (
  .F(lut_f_1992),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1992.INIT = 16'h8000;
LUT4 lut_inst_1993 (
  .F(lut_f_1993),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1993.INIT = 16'h8000;
LUT4 lut_inst_1994 (
  .F(lut_f_1994),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1994.INIT = 16'h8000;
LUT4 lut_inst_1995 (
  .F(lut_f_1995),
  .I0(lut_f_1992),
  .I1(lut_f_1993),
  .I2(lut_f_1994),
  .I3(gw_vcc)
);
defparam lut_inst_1995.INIT = 16'h8000;
LUT4 lut_inst_1996 (
  .F(lut_f_1996),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_1996.INIT = 16'h8000;
LUT4 lut_inst_1997 (
  .F(lut_f_1997),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_1997.INIT = 16'h8000;
LUT4 lut_inst_1998 (
  .F(lut_f_1998),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1998.INIT = 16'h8000;
LUT4 lut_inst_1999 (
  .F(lut_f_1999),
  .I0(lut_f_1996),
  .I1(lut_f_1997),
  .I2(lut_f_1998),
  .I3(gw_vcc)
);
defparam lut_inst_1999.INIT = 16'h8000;
LUT4 lut_inst_2000 (
  .F(lut_f_2000),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2000.INIT = 16'h8000;
LUT4 lut_inst_2001 (
  .F(lut_f_2001),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2001.INIT = 16'h8000;
LUT4 lut_inst_2002 (
  .F(lut_f_2002),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_2002.INIT = 16'h8000;
LUT4 lut_inst_2003 (
  .F(lut_f_2003),
  .I0(lut_f_2000),
  .I1(lut_f_2001),
  .I2(lut_f_2002),
  .I3(gw_vcc)
);
defparam lut_inst_2003.INIT = 16'h8000;
LUT4 lut_inst_2004 (
  .F(lut_f_2004),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2004.INIT = 16'h8000;
LUT4 lut_inst_2005 (
  .F(lut_f_2005),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2005.INIT = 16'h8000;
LUT4 lut_inst_2006 (
  .F(lut_f_2006),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_2006.INIT = 16'h8000;
LUT4 lut_inst_2007 (
  .F(lut_f_2007),
  .I0(lut_f_2004),
  .I1(lut_f_2005),
  .I2(lut_f_2006),
  .I3(gw_vcc)
);
defparam lut_inst_2007.INIT = 16'h8000;
LUT4 lut_inst_2008 (
  .F(lut_f_2008),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2008.INIT = 16'h8000;
LUT4 lut_inst_2009 (
  .F(lut_f_2009),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2009.INIT = 16'h8000;
LUT4 lut_inst_2010 (
  .F(lut_f_2010),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_2010.INIT = 16'h8000;
LUT4 lut_inst_2011 (
  .F(lut_f_2011),
  .I0(lut_f_2008),
  .I1(lut_f_2009),
  .I2(lut_f_2010),
  .I3(gw_vcc)
);
defparam lut_inst_2011.INIT = 16'h8000;
LUT4 lut_inst_2012 (
  .F(lut_f_2012),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2012.INIT = 16'h8000;
LUT4 lut_inst_2013 (
  .F(lut_f_2013),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2013.INIT = 16'h8000;
LUT4 lut_inst_2014 (
  .F(lut_f_2014),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_2014.INIT = 16'h8000;
LUT4 lut_inst_2015 (
  .F(lut_f_2015),
  .I0(lut_f_2012),
  .I1(lut_f_2013),
  .I2(lut_f_2014),
  .I3(gw_vcc)
);
defparam lut_inst_2015.INIT = 16'h8000;
LUT4 lut_inst_2016 (
  .F(lut_f_2016),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2016.INIT = 16'h8000;
LUT4 lut_inst_2017 (
  .F(lut_f_2017),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2017.INIT = 16'h8000;
LUT4 lut_inst_2018 (
  .F(lut_f_2018),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_2018.INIT = 16'h8000;
LUT4 lut_inst_2019 (
  .F(lut_f_2019),
  .I0(lut_f_2016),
  .I1(lut_f_2017),
  .I2(lut_f_2018),
  .I3(gw_vcc)
);
defparam lut_inst_2019.INIT = 16'h8000;
LUT4 lut_inst_2020 (
  .F(lut_f_2020),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2020.INIT = 16'h8000;
LUT4 lut_inst_2021 (
  .F(lut_f_2021),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2021.INIT = 16'h8000;
LUT4 lut_inst_2022 (
  .F(lut_f_2022),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_2022.INIT = 16'h8000;
LUT4 lut_inst_2023 (
  .F(lut_f_2023),
  .I0(lut_f_2020),
  .I1(lut_f_2021),
  .I2(lut_f_2022),
  .I3(gw_vcc)
);
defparam lut_inst_2023.INIT = 16'h8000;
LUT4 lut_inst_2024 (
  .F(lut_f_2024),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2024.INIT = 16'h8000;
LUT4 lut_inst_2025 (
  .F(lut_f_2025),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2025.INIT = 16'h8000;
LUT4 lut_inst_2026 (
  .F(lut_f_2026),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_2026.INIT = 16'h8000;
LUT4 lut_inst_2027 (
  .F(lut_f_2027),
  .I0(lut_f_2024),
  .I1(lut_f_2025),
  .I2(lut_f_2026),
  .I3(gw_vcc)
);
defparam lut_inst_2027.INIT = 16'h8000;
LUT4 lut_inst_2028 (
  .F(lut_f_2028),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2028.INIT = 16'h8000;
LUT4 lut_inst_2029 (
  .F(lut_f_2029),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2029.INIT = 16'h8000;
LUT4 lut_inst_2030 (
  .F(lut_f_2030),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_2030.INIT = 16'h8000;
LUT4 lut_inst_2031 (
  .F(lut_f_2031),
  .I0(lut_f_2028),
  .I1(lut_f_2029),
  .I2(lut_f_2030),
  .I3(gw_vcc)
);
defparam lut_inst_2031.INIT = 16'h8000;
LUT4 lut_inst_2032 (
  .F(lut_f_2032),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2032.INIT = 16'h8000;
LUT4 lut_inst_2033 (
  .F(lut_f_2033),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2033.INIT = 16'h8000;
LUT4 lut_inst_2034 (
  .F(lut_f_2034),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_2034.INIT = 16'h8000;
LUT4 lut_inst_2035 (
  .F(lut_f_2035),
  .I0(lut_f_2032),
  .I1(lut_f_2033),
  .I2(lut_f_2034),
  .I3(gw_vcc)
);
defparam lut_inst_2035.INIT = 16'h8000;
LUT4 lut_inst_2036 (
  .F(lut_f_2036),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2036.INIT = 16'h8000;
LUT4 lut_inst_2037 (
  .F(lut_f_2037),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2037.INIT = 16'h8000;
LUT4 lut_inst_2038 (
  .F(lut_f_2038),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_2038.INIT = 16'h8000;
LUT4 lut_inst_2039 (
  .F(lut_f_2039),
  .I0(lut_f_2036),
  .I1(lut_f_2037),
  .I2(lut_f_2038),
  .I3(gw_vcc)
);
defparam lut_inst_2039.INIT = 16'h8000;
LUT4 lut_inst_2040 (
  .F(lut_f_2040),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2040.INIT = 16'h8000;
LUT4 lut_inst_2041 (
  .F(lut_f_2041),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2041.INIT = 16'h8000;
LUT4 lut_inst_2042 (
  .F(lut_f_2042),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_2042.INIT = 16'h8000;
LUT4 lut_inst_2043 (
  .F(lut_f_2043),
  .I0(lut_f_2040),
  .I1(lut_f_2041),
  .I2(lut_f_2042),
  .I3(gw_vcc)
);
defparam lut_inst_2043.INIT = 16'h8000;
LUT4 lut_inst_2044 (
  .F(lut_f_2044),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2044.INIT = 16'h8000;
LUT4 lut_inst_2045 (
  .F(lut_f_2045),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2045.INIT = 16'h8000;
LUT4 lut_inst_2046 (
  .F(lut_f_2046),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad13_inv),
  .I3(gw_vcc)
);
defparam lut_inst_2046.INIT = 16'h8000;
LUT4 lut_inst_2047 (
  .F(lut_f_2047),
  .I0(lut_f_2044),
  .I1(lut_f_2045),
  .I2(lut_f_2046),
  .I3(gw_vcc)
);
defparam lut_inst_2047.INIT = 16'h8000;
LUT4 lut_inst_2048 (
  .F(lut_f_2048),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2048.INIT = 16'h8000;
LUT4 lut_inst_2049 (
  .F(lut_f_2049),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2049.INIT = 16'h8000;
LUT4 lut_inst_2050 (
  .F(lut_f_2050),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2050.INIT = 16'h8000;
LUT4 lut_inst_2051 (
  .F(lut_f_2051),
  .I0(lut_f_2048),
  .I1(lut_f_2049),
  .I2(lut_f_2050),
  .I3(gw_vcc)
);
defparam lut_inst_2051.INIT = 16'h8000;
LUT4 lut_inst_2052 (
  .F(lut_f_2052),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2052.INIT = 16'h8000;
LUT4 lut_inst_2053 (
  .F(lut_f_2053),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2053.INIT = 16'h8000;
LUT4 lut_inst_2054 (
  .F(lut_f_2054),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2054.INIT = 16'h8000;
LUT4 lut_inst_2055 (
  .F(lut_f_2055),
  .I0(lut_f_2052),
  .I1(lut_f_2053),
  .I2(lut_f_2054),
  .I3(gw_vcc)
);
defparam lut_inst_2055.INIT = 16'h8000;
LUT4 lut_inst_2056 (
  .F(lut_f_2056),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2056.INIT = 16'h8000;
LUT4 lut_inst_2057 (
  .F(lut_f_2057),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2057.INIT = 16'h8000;
LUT4 lut_inst_2058 (
  .F(lut_f_2058),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2058.INIT = 16'h8000;
LUT4 lut_inst_2059 (
  .F(lut_f_2059),
  .I0(lut_f_2056),
  .I1(lut_f_2057),
  .I2(lut_f_2058),
  .I3(gw_vcc)
);
defparam lut_inst_2059.INIT = 16'h8000;
LUT4 lut_inst_2060 (
  .F(lut_f_2060),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2060.INIT = 16'h8000;
LUT4 lut_inst_2061 (
  .F(lut_f_2061),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2061.INIT = 16'h8000;
LUT4 lut_inst_2062 (
  .F(lut_f_2062),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2062.INIT = 16'h8000;
LUT4 lut_inst_2063 (
  .F(lut_f_2063),
  .I0(lut_f_2060),
  .I1(lut_f_2061),
  .I2(lut_f_2062),
  .I3(gw_vcc)
);
defparam lut_inst_2063.INIT = 16'h8000;
LUT4 lut_inst_2064 (
  .F(lut_f_2064),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2064.INIT = 16'h8000;
LUT4 lut_inst_2065 (
  .F(lut_f_2065),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2065.INIT = 16'h8000;
LUT4 lut_inst_2066 (
  .F(lut_f_2066),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2066.INIT = 16'h8000;
LUT4 lut_inst_2067 (
  .F(lut_f_2067),
  .I0(lut_f_2064),
  .I1(lut_f_2065),
  .I2(lut_f_2066),
  .I3(gw_vcc)
);
defparam lut_inst_2067.INIT = 16'h8000;
LUT4 lut_inst_2068 (
  .F(lut_f_2068),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2068.INIT = 16'h8000;
LUT4 lut_inst_2069 (
  .F(lut_f_2069),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2069.INIT = 16'h8000;
LUT4 lut_inst_2070 (
  .F(lut_f_2070),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2070.INIT = 16'h8000;
LUT4 lut_inst_2071 (
  .F(lut_f_2071),
  .I0(lut_f_2068),
  .I1(lut_f_2069),
  .I2(lut_f_2070),
  .I3(gw_vcc)
);
defparam lut_inst_2071.INIT = 16'h8000;
LUT4 lut_inst_2072 (
  .F(lut_f_2072),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2072.INIT = 16'h8000;
LUT4 lut_inst_2073 (
  .F(lut_f_2073),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2073.INIT = 16'h8000;
LUT4 lut_inst_2074 (
  .F(lut_f_2074),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2074.INIT = 16'h8000;
LUT4 lut_inst_2075 (
  .F(lut_f_2075),
  .I0(lut_f_2072),
  .I1(lut_f_2073),
  .I2(lut_f_2074),
  .I3(gw_vcc)
);
defparam lut_inst_2075.INIT = 16'h8000;
LUT4 lut_inst_2076 (
  .F(lut_f_2076),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2076.INIT = 16'h8000;
LUT4 lut_inst_2077 (
  .F(lut_f_2077),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2077.INIT = 16'h8000;
LUT4 lut_inst_2078 (
  .F(lut_f_2078),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2078.INIT = 16'h8000;
LUT4 lut_inst_2079 (
  .F(lut_f_2079),
  .I0(lut_f_2076),
  .I1(lut_f_2077),
  .I2(lut_f_2078),
  .I3(gw_vcc)
);
defparam lut_inst_2079.INIT = 16'h8000;
LUT4 lut_inst_2080 (
  .F(lut_f_2080),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2080.INIT = 16'h8000;
LUT4 lut_inst_2081 (
  .F(lut_f_2081),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2081.INIT = 16'h8000;
LUT4 lut_inst_2082 (
  .F(lut_f_2082),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2082.INIT = 16'h8000;
LUT4 lut_inst_2083 (
  .F(lut_f_2083),
  .I0(lut_f_2080),
  .I1(lut_f_2081),
  .I2(lut_f_2082),
  .I3(gw_vcc)
);
defparam lut_inst_2083.INIT = 16'h8000;
LUT4 lut_inst_2084 (
  .F(lut_f_2084),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2084.INIT = 16'h8000;
LUT4 lut_inst_2085 (
  .F(lut_f_2085),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2085.INIT = 16'h8000;
LUT4 lut_inst_2086 (
  .F(lut_f_2086),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2086.INIT = 16'h8000;
LUT4 lut_inst_2087 (
  .F(lut_f_2087),
  .I0(lut_f_2084),
  .I1(lut_f_2085),
  .I2(lut_f_2086),
  .I3(gw_vcc)
);
defparam lut_inst_2087.INIT = 16'h8000;
LUT4 lut_inst_2088 (
  .F(lut_f_2088),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2088.INIT = 16'h8000;
LUT4 lut_inst_2089 (
  .F(lut_f_2089),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2089.INIT = 16'h8000;
LUT4 lut_inst_2090 (
  .F(lut_f_2090),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2090.INIT = 16'h8000;
LUT4 lut_inst_2091 (
  .F(lut_f_2091),
  .I0(lut_f_2088),
  .I1(lut_f_2089),
  .I2(lut_f_2090),
  .I3(gw_vcc)
);
defparam lut_inst_2091.INIT = 16'h8000;
LUT4 lut_inst_2092 (
  .F(lut_f_2092),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2092.INIT = 16'h8000;
LUT4 lut_inst_2093 (
  .F(lut_f_2093),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2093.INIT = 16'h8000;
LUT4 lut_inst_2094 (
  .F(lut_f_2094),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2094.INIT = 16'h8000;
LUT4 lut_inst_2095 (
  .F(lut_f_2095),
  .I0(lut_f_2092),
  .I1(lut_f_2093),
  .I2(lut_f_2094),
  .I3(gw_vcc)
);
defparam lut_inst_2095.INIT = 16'h8000;
LUT4 lut_inst_2096 (
  .F(lut_f_2096),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2096.INIT = 16'h8000;
LUT4 lut_inst_2097 (
  .F(lut_f_2097),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2097.INIT = 16'h8000;
LUT4 lut_inst_2098 (
  .F(lut_f_2098),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2098.INIT = 16'h8000;
LUT4 lut_inst_2099 (
  .F(lut_f_2099),
  .I0(lut_f_2096),
  .I1(lut_f_2097),
  .I2(lut_f_2098),
  .I3(gw_vcc)
);
defparam lut_inst_2099.INIT = 16'h8000;
LUT4 lut_inst_2100 (
  .F(lut_f_2100),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2100.INIT = 16'h8000;
LUT4 lut_inst_2101 (
  .F(lut_f_2101),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2101.INIT = 16'h8000;
LUT4 lut_inst_2102 (
  .F(lut_f_2102),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2102.INIT = 16'h8000;
LUT4 lut_inst_2103 (
  .F(lut_f_2103),
  .I0(lut_f_2100),
  .I1(lut_f_2101),
  .I2(lut_f_2102),
  .I3(gw_vcc)
);
defparam lut_inst_2103.INIT = 16'h8000;
LUT4 lut_inst_2104 (
  .F(lut_f_2104),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2104.INIT = 16'h8000;
LUT4 lut_inst_2105 (
  .F(lut_f_2105),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2105.INIT = 16'h8000;
LUT4 lut_inst_2106 (
  .F(lut_f_2106),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2106.INIT = 16'h8000;
LUT4 lut_inst_2107 (
  .F(lut_f_2107),
  .I0(lut_f_2104),
  .I1(lut_f_2105),
  .I2(lut_f_2106),
  .I3(gw_vcc)
);
defparam lut_inst_2107.INIT = 16'h8000;
LUT4 lut_inst_2108 (
  .F(lut_f_2108),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2108.INIT = 16'h8000;
LUT4 lut_inst_2109 (
  .F(lut_f_2109),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2109.INIT = 16'h8000;
LUT4 lut_inst_2110 (
  .F(lut_f_2110),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2110.INIT = 16'h8000;
LUT4 lut_inst_2111 (
  .F(lut_f_2111),
  .I0(lut_f_2108),
  .I1(lut_f_2109),
  .I2(lut_f_2110),
  .I3(gw_vcc)
);
defparam lut_inst_2111.INIT = 16'h8000;
LUT4 lut_inst_2112 (
  .F(lut_f_2112),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2112.INIT = 16'h8000;
LUT4 lut_inst_2113 (
  .F(lut_f_2113),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2113.INIT = 16'h8000;
LUT4 lut_inst_2114 (
  .F(lut_f_2114),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2114.INIT = 16'h8000;
LUT4 lut_inst_2115 (
  .F(lut_f_2115),
  .I0(lut_f_2112),
  .I1(lut_f_2113),
  .I2(lut_f_2114),
  .I3(gw_vcc)
);
defparam lut_inst_2115.INIT = 16'h8000;
LUT4 lut_inst_2116 (
  .F(lut_f_2116),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2116.INIT = 16'h8000;
LUT4 lut_inst_2117 (
  .F(lut_f_2117),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2117.INIT = 16'h8000;
LUT4 lut_inst_2118 (
  .F(lut_f_2118),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2118.INIT = 16'h8000;
LUT4 lut_inst_2119 (
  .F(lut_f_2119),
  .I0(lut_f_2116),
  .I1(lut_f_2117),
  .I2(lut_f_2118),
  .I3(gw_vcc)
);
defparam lut_inst_2119.INIT = 16'h8000;
LUT4 lut_inst_2120 (
  .F(lut_f_2120),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2120.INIT = 16'h8000;
LUT4 lut_inst_2121 (
  .F(lut_f_2121),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2121.INIT = 16'h8000;
LUT4 lut_inst_2122 (
  .F(lut_f_2122),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2122.INIT = 16'h8000;
LUT4 lut_inst_2123 (
  .F(lut_f_2123),
  .I0(lut_f_2120),
  .I1(lut_f_2121),
  .I2(lut_f_2122),
  .I3(gw_vcc)
);
defparam lut_inst_2123.INIT = 16'h8000;
LUT4 lut_inst_2124 (
  .F(lut_f_2124),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2124.INIT = 16'h8000;
LUT4 lut_inst_2125 (
  .F(lut_f_2125),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2125.INIT = 16'h8000;
LUT4 lut_inst_2126 (
  .F(lut_f_2126),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2126.INIT = 16'h8000;
LUT4 lut_inst_2127 (
  .F(lut_f_2127),
  .I0(lut_f_2124),
  .I1(lut_f_2125),
  .I2(lut_f_2126),
  .I3(gw_vcc)
);
defparam lut_inst_2127.INIT = 16'h8000;
LUT4 lut_inst_2128 (
  .F(lut_f_2128),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2128.INIT = 16'h8000;
LUT4 lut_inst_2129 (
  .F(lut_f_2129),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2129.INIT = 16'h8000;
LUT4 lut_inst_2130 (
  .F(lut_f_2130),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2130.INIT = 16'h8000;
LUT4 lut_inst_2131 (
  .F(lut_f_2131),
  .I0(lut_f_2128),
  .I1(lut_f_2129),
  .I2(lut_f_2130),
  .I3(gw_vcc)
);
defparam lut_inst_2131.INIT = 16'h8000;
LUT4 lut_inst_2132 (
  .F(lut_f_2132),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2132.INIT = 16'h8000;
LUT4 lut_inst_2133 (
  .F(lut_f_2133),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2133.INIT = 16'h8000;
LUT4 lut_inst_2134 (
  .F(lut_f_2134),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2134.INIT = 16'h8000;
LUT4 lut_inst_2135 (
  .F(lut_f_2135),
  .I0(lut_f_2132),
  .I1(lut_f_2133),
  .I2(lut_f_2134),
  .I3(gw_vcc)
);
defparam lut_inst_2135.INIT = 16'h8000;
LUT4 lut_inst_2136 (
  .F(lut_f_2136),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2136.INIT = 16'h8000;
LUT4 lut_inst_2137 (
  .F(lut_f_2137),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2137.INIT = 16'h8000;
LUT4 lut_inst_2138 (
  .F(lut_f_2138),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2138.INIT = 16'h8000;
LUT4 lut_inst_2139 (
  .F(lut_f_2139),
  .I0(lut_f_2136),
  .I1(lut_f_2137),
  .I2(lut_f_2138),
  .I3(gw_vcc)
);
defparam lut_inst_2139.INIT = 16'h8000;
LUT4 lut_inst_2140 (
  .F(lut_f_2140),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2140.INIT = 16'h8000;
LUT4 lut_inst_2141 (
  .F(lut_f_2141),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2141.INIT = 16'h8000;
LUT4 lut_inst_2142 (
  .F(lut_f_2142),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2142.INIT = 16'h8000;
LUT4 lut_inst_2143 (
  .F(lut_f_2143),
  .I0(lut_f_2140),
  .I1(lut_f_2141),
  .I2(lut_f_2142),
  .I3(gw_vcc)
);
defparam lut_inst_2143.INIT = 16'h8000;
LUT4 lut_inst_2144 (
  .F(lut_f_2144),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2144.INIT = 16'h8000;
LUT4 lut_inst_2145 (
  .F(lut_f_2145),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2145.INIT = 16'h8000;
LUT4 lut_inst_2146 (
  .F(lut_f_2146),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2146.INIT = 16'h8000;
LUT4 lut_inst_2147 (
  .F(lut_f_2147),
  .I0(lut_f_2144),
  .I1(lut_f_2145),
  .I2(lut_f_2146),
  .I3(gw_vcc)
);
defparam lut_inst_2147.INIT = 16'h8000;
LUT4 lut_inst_2148 (
  .F(lut_f_2148),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2148.INIT = 16'h8000;
LUT4 lut_inst_2149 (
  .F(lut_f_2149),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2149.INIT = 16'h8000;
LUT4 lut_inst_2150 (
  .F(lut_f_2150),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2150.INIT = 16'h8000;
LUT4 lut_inst_2151 (
  .F(lut_f_2151),
  .I0(lut_f_2148),
  .I1(lut_f_2149),
  .I2(lut_f_2150),
  .I3(gw_vcc)
);
defparam lut_inst_2151.INIT = 16'h8000;
LUT4 lut_inst_2152 (
  .F(lut_f_2152),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2152.INIT = 16'h8000;
LUT4 lut_inst_2153 (
  .F(lut_f_2153),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2153.INIT = 16'h8000;
LUT4 lut_inst_2154 (
  .F(lut_f_2154),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2154.INIT = 16'h8000;
LUT4 lut_inst_2155 (
  .F(lut_f_2155),
  .I0(lut_f_2152),
  .I1(lut_f_2153),
  .I2(lut_f_2154),
  .I3(gw_vcc)
);
defparam lut_inst_2155.INIT = 16'h8000;
LUT4 lut_inst_2156 (
  .F(lut_f_2156),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2156.INIT = 16'h8000;
LUT4 lut_inst_2157 (
  .F(lut_f_2157),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2157.INIT = 16'h8000;
LUT4 lut_inst_2158 (
  .F(lut_f_2158),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2158.INIT = 16'h8000;
LUT4 lut_inst_2159 (
  .F(lut_f_2159),
  .I0(lut_f_2156),
  .I1(lut_f_2157),
  .I2(lut_f_2158),
  .I3(gw_vcc)
);
defparam lut_inst_2159.INIT = 16'h8000;
LUT4 lut_inst_2160 (
  .F(lut_f_2160),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2160.INIT = 16'h8000;
LUT4 lut_inst_2161 (
  .F(lut_f_2161),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2161.INIT = 16'h8000;
LUT4 lut_inst_2162 (
  .F(lut_f_2162),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2162.INIT = 16'h8000;
LUT4 lut_inst_2163 (
  .F(lut_f_2163),
  .I0(lut_f_2160),
  .I1(lut_f_2161),
  .I2(lut_f_2162),
  .I3(gw_vcc)
);
defparam lut_inst_2163.INIT = 16'h8000;
LUT4 lut_inst_2164 (
  .F(lut_f_2164),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2164.INIT = 16'h8000;
LUT4 lut_inst_2165 (
  .F(lut_f_2165),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2165.INIT = 16'h8000;
LUT4 lut_inst_2166 (
  .F(lut_f_2166),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2166.INIT = 16'h8000;
LUT4 lut_inst_2167 (
  .F(lut_f_2167),
  .I0(lut_f_2164),
  .I1(lut_f_2165),
  .I2(lut_f_2166),
  .I3(gw_vcc)
);
defparam lut_inst_2167.INIT = 16'h8000;
LUT4 lut_inst_2168 (
  .F(lut_f_2168),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2168.INIT = 16'h8000;
LUT4 lut_inst_2169 (
  .F(lut_f_2169),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2169.INIT = 16'h8000;
LUT4 lut_inst_2170 (
  .F(lut_f_2170),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2170.INIT = 16'h8000;
LUT4 lut_inst_2171 (
  .F(lut_f_2171),
  .I0(lut_f_2168),
  .I1(lut_f_2169),
  .I2(lut_f_2170),
  .I3(gw_vcc)
);
defparam lut_inst_2171.INIT = 16'h8000;
LUT4 lut_inst_2172 (
  .F(lut_f_2172),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2172.INIT = 16'h8000;
LUT4 lut_inst_2173 (
  .F(lut_f_2173),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2173.INIT = 16'h8000;
LUT4 lut_inst_2174 (
  .F(lut_f_2174),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2174.INIT = 16'h8000;
LUT4 lut_inst_2175 (
  .F(lut_f_2175),
  .I0(lut_f_2172),
  .I1(lut_f_2173),
  .I2(lut_f_2174),
  .I3(gw_vcc)
);
defparam lut_inst_2175.INIT = 16'h8000;
LUT4 lut_inst_2176 (
  .F(lut_f_2176),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2176.INIT = 16'h8000;
LUT4 lut_inst_2177 (
  .F(lut_f_2177),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2177.INIT = 16'h8000;
LUT4 lut_inst_2178 (
  .F(lut_f_2178),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2178.INIT = 16'h8000;
LUT4 lut_inst_2179 (
  .F(lut_f_2179),
  .I0(lut_f_2176),
  .I1(lut_f_2177),
  .I2(lut_f_2178),
  .I3(gw_vcc)
);
defparam lut_inst_2179.INIT = 16'h8000;
LUT4 lut_inst_2180 (
  .F(lut_f_2180),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2180.INIT = 16'h8000;
LUT4 lut_inst_2181 (
  .F(lut_f_2181),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2181.INIT = 16'h8000;
LUT4 lut_inst_2182 (
  .F(lut_f_2182),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2182.INIT = 16'h8000;
LUT4 lut_inst_2183 (
  .F(lut_f_2183),
  .I0(lut_f_2180),
  .I1(lut_f_2181),
  .I2(lut_f_2182),
  .I3(gw_vcc)
);
defparam lut_inst_2183.INIT = 16'h8000;
LUT4 lut_inst_2184 (
  .F(lut_f_2184),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2184.INIT = 16'h8000;
LUT4 lut_inst_2185 (
  .F(lut_f_2185),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2185.INIT = 16'h8000;
LUT4 lut_inst_2186 (
  .F(lut_f_2186),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2186.INIT = 16'h8000;
LUT4 lut_inst_2187 (
  .F(lut_f_2187),
  .I0(lut_f_2184),
  .I1(lut_f_2185),
  .I2(lut_f_2186),
  .I3(gw_vcc)
);
defparam lut_inst_2187.INIT = 16'h8000;
LUT4 lut_inst_2188 (
  .F(lut_f_2188),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2188.INIT = 16'h8000;
LUT4 lut_inst_2189 (
  .F(lut_f_2189),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2189.INIT = 16'h8000;
LUT4 lut_inst_2190 (
  .F(lut_f_2190),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2190.INIT = 16'h8000;
LUT4 lut_inst_2191 (
  .F(lut_f_2191),
  .I0(lut_f_2188),
  .I1(lut_f_2189),
  .I2(lut_f_2190),
  .I3(gw_vcc)
);
defparam lut_inst_2191.INIT = 16'h8000;
LUT4 lut_inst_2192 (
  .F(lut_f_2192),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2192.INIT = 16'h8000;
LUT4 lut_inst_2193 (
  .F(lut_f_2193),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2193.INIT = 16'h8000;
LUT4 lut_inst_2194 (
  .F(lut_f_2194),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2194.INIT = 16'h8000;
LUT4 lut_inst_2195 (
  .F(lut_f_2195),
  .I0(lut_f_2192),
  .I1(lut_f_2193),
  .I2(lut_f_2194),
  .I3(gw_vcc)
);
defparam lut_inst_2195.INIT = 16'h8000;
LUT4 lut_inst_2196 (
  .F(lut_f_2196),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2196.INIT = 16'h8000;
LUT4 lut_inst_2197 (
  .F(lut_f_2197),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2197.INIT = 16'h8000;
LUT4 lut_inst_2198 (
  .F(lut_f_2198),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2198.INIT = 16'h8000;
LUT4 lut_inst_2199 (
  .F(lut_f_2199),
  .I0(lut_f_2196),
  .I1(lut_f_2197),
  .I2(lut_f_2198),
  .I3(gw_vcc)
);
defparam lut_inst_2199.INIT = 16'h8000;
LUT4 lut_inst_2200 (
  .F(lut_f_2200),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2200.INIT = 16'h8000;
LUT4 lut_inst_2201 (
  .F(lut_f_2201),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2201.INIT = 16'h8000;
LUT4 lut_inst_2202 (
  .F(lut_f_2202),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2202.INIT = 16'h8000;
LUT4 lut_inst_2203 (
  .F(lut_f_2203),
  .I0(lut_f_2200),
  .I1(lut_f_2201),
  .I2(lut_f_2202),
  .I3(gw_vcc)
);
defparam lut_inst_2203.INIT = 16'h8000;
LUT4 lut_inst_2204 (
  .F(lut_f_2204),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2204.INIT = 16'h8000;
LUT4 lut_inst_2205 (
  .F(lut_f_2205),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2205.INIT = 16'h8000;
LUT4 lut_inst_2206 (
  .F(lut_f_2206),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2206.INIT = 16'h8000;
LUT4 lut_inst_2207 (
  .F(lut_f_2207),
  .I0(lut_f_2204),
  .I1(lut_f_2205),
  .I2(lut_f_2206),
  .I3(gw_vcc)
);
defparam lut_inst_2207.INIT = 16'h8000;
LUT4 lut_inst_2208 (
  .F(lut_f_2208),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2208.INIT = 16'h8000;
LUT4 lut_inst_2209 (
  .F(lut_f_2209),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2209.INIT = 16'h8000;
LUT4 lut_inst_2210 (
  .F(lut_f_2210),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2210.INIT = 16'h8000;
LUT4 lut_inst_2211 (
  .F(lut_f_2211),
  .I0(lut_f_2208),
  .I1(lut_f_2209),
  .I2(lut_f_2210),
  .I3(gw_vcc)
);
defparam lut_inst_2211.INIT = 16'h8000;
LUT4 lut_inst_2212 (
  .F(lut_f_2212),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2212.INIT = 16'h8000;
LUT4 lut_inst_2213 (
  .F(lut_f_2213),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2213.INIT = 16'h8000;
LUT4 lut_inst_2214 (
  .F(lut_f_2214),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2214.INIT = 16'h8000;
LUT4 lut_inst_2215 (
  .F(lut_f_2215),
  .I0(lut_f_2212),
  .I1(lut_f_2213),
  .I2(lut_f_2214),
  .I3(gw_vcc)
);
defparam lut_inst_2215.INIT = 16'h8000;
LUT4 lut_inst_2216 (
  .F(lut_f_2216),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2216.INIT = 16'h8000;
LUT4 lut_inst_2217 (
  .F(lut_f_2217),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2217.INIT = 16'h8000;
LUT4 lut_inst_2218 (
  .F(lut_f_2218),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2218.INIT = 16'h8000;
LUT4 lut_inst_2219 (
  .F(lut_f_2219),
  .I0(lut_f_2216),
  .I1(lut_f_2217),
  .I2(lut_f_2218),
  .I3(gw_vcc)
);
defparam lut_inst_2219.INIT = 16'h8000;
LUT4 lut_inst_2220 (
  .F(lut_f_2220),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2220.INIT = 16'h8000;
LUT4 lut_inst_2221 (
  .F(lut_f_2221),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2221.INIT = 16'h8000;
LUT4 lut_inst_2222 (
  .F(lut_f_2222),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2222.INIT = 16'h8000;
LUT4 lut_inst_2223 (
  .F(lut_f_2223),
  .I0(lut_f_2220),
  .I1(lut_f_2221),
  .I2(lut_f_2222),
  .I3(gw_vcc)
);
defparam lut_inst_2223.INIT = 16'h8000;
LUT4 lut_inst_2224 (
  .F(lut_f_2224),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2224.INIT = 16'h8000;
LUT4 lut_inst_2225 (
  .F(lut_f_2225),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2225.INIT = 16'h8000;
LUT4 lut_inst_2226 (
  .F(lut_f_2226),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2226.INIT = 16'h8000;
LUT4 lut_inst_2227 (
  .F(lut_f_2227),
  .I0(lut_f_2224),
  .I1(lut_f_2225),
  .I2(lut_f_2226),
  .I3(gw_vcc)
);
defparam lut_inst_2227.INIT = 16'h8000;
LUT4 lut_inst_2228 (
  .F(lut_f_2228),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2228.INIT = 16'h8000;
LUT4 lut_inst_2229 (
  .F(lut_f_2229),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2229.INIT = 16'h8000;
LUT4 lut_inst_2230 (
  .F(lut_f_2230),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2230.INIT = 16'h8000;
LUT4 lut_inst_2231 (
  .F(lut_f_2231),
  .I0(lut_f_2228),
  .I1(lut_f_2229),
  .I2(lut_f_2230),
  .I3(gw_vcc)
);
defparam lut_inst_2231.INIT = 16'h8000;
LUT4 lut_inst_2232 (
  .F(lut_f_2232),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2232.INIT = 16'h8000;
LUT4 lut_inst_2233 (
  .F(lut_f_2233),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2233.INIT = 16'h8000;
LUT4 lut_inst_2234 (
  .F(lut_f_2234),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2234.INIT = 16'h8000;
LUT4 lut_inst_2235 (
  .F(lut_f_2235),
  .I0(lut_f_2232),
  .I1(lut_f_2233),
  .I2(lut_f_2234),
  .I3(gw_vcc)
);
defparam lut_inst_2235.INIT = 16'h8000;
LUT4 lut_inst_2236 (
  .F(lut_f_2236),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2236.INIT = 16'h8000;
LUT4 lut_inst_2237 (
  .F(lut_f_2237),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2237.INIT = 16'h8000;
LUT4 lut_inst_2238 (
  .F(lut_f_2238),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2238.INIT = 16'h8000;
LUT4 lut_inst_2239 (
  .F(lut_f_2239),
  .I0(lut_f_2236),
  .I1(lut_f_2237),
  .I2(lut_f_2238),
  .I3(gw_vcc)
);
defparam lut_inst_2239.INIT = 16'h8000;
LUT4 lut_inst_2240 (
  .F(lut_f_2240),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2240.INIT = 16'h8000;
LUT4 lut_inst_2241 (
  .F(lut_f_2241),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2241.INIT = 16'h8000;
LUT4 lut_inst_2242 (
  .F(lut_f_2242),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2242.INIT = 16'h8000;
LUT4 lut_inst_2243 (
  .F(lut_f_2243),
  .I0(lut_f_2240),
  .I1(lut_f_2241),
  .I2(lut_f_2242),
  .I3(gw_vcc)
);
defparam lut_inst_2243.INIT = 16'h8000;
LUT4 lut_inst_2244 (
  .F(lut_f_2244),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2244.INIT = 16'h8000;
LUT4 lut_inst_2245 (
  .F(lut_f_2245),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2245.INIT = 16'h8000;
LUT4 lut_inst_2246 (
  .F(lut_f_2246),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2246.INIT = 16'h8000;
LUT4 lut_inst_2247 (
  .F(lut_f_2247),
  .I0(lut_f_2244),
  .I1(lut_f_2245),
  .I2(lut_f_2246),
  .I3(gw_vcc)
);
defparam lut_inst_2247.INIT = 16'h8000;
LUT4 lut_inst_2248 (
  .F(lut_f_2248),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2248.INIT = 16'h8000;
LUT4 lut_inst_2249 (
  .F(lut_f_2249),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2249.INIT = 16'h8000;
LUT4 lut_inst_2250 (
  .F(lut_f_2250),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2250.INIT = 16'h8000;
LUT4 lut_inst_2251 (
  .F(lut_f_2251),
  .I0(lut_f_2248),
  .I1(lut_f_2249),
  .I2(lut_f_2250),
  .I3(gw_vcc)
);
defparam lut_inst_2251.INIT = 16'h8000;
LUT4 lut_inst_2252 (
  .F(lut_f_2252),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2252.INIT = 16'h8000;
LUT4 lut_inst_2253 (
  .F(lut_f_2253),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2253.INIT = 16'h8000;
LUT4 lut_inst_2254 (
  .F(lut_f_2254),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2254.INIT = 16'h8000;
LUT4 lut_inst_2255 (
  .F(lut_f_2255),
  .I0(lut_f_2252),
  .I1(lut_f_2253),
  .I2(lut_f_2254),
  .I3(gw_vcc)
);
defparam lut_inst_2255.INIT = 16'h8000;
LUT4 lut_inst_2256 (
  .F(lut_f_2256),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2256.INIT = 16'h8000;
LUT4 lut_inst_2257 (
  .F(lut_f_2257),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2257.INIT = 16'h8000;
LUT4 lut_inst_2258 (
  .F(lut_f_2258),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2258.INIT = 16'h8000;
LUT4 lut_inst_2259 (
  .F(lut_f_2259),
  .I0(lut_f_2256),
  .I1(lut_f_2257),
  .I2(lut_f_2258),
  .I3(gw_vcc)
);
defparam lut_inst_2259.INIT = 16'h8000;
LUT4 lut_inst_2260 (
  .F(lut_f_2260),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2260.INIT = 16'h8000;
LUT4 lut_inst_2261 (
  .F(lut_f_2261),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2261.INIT = 16'h8000;
LUT4 lut_inst_2262 (
  .F(lut_f_2262),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2262.INIT = 16'h8000;
LUT4 lut_inst_2263 (
  .F(lut_f_2263),
  .I0(lut_f_2260),
  .I1(lut_f_2261),
  .I2(lut_f_2262),
  .I3(gw_vcc)
);
defparam lut_inst_2263.INIT = 16'h8000;
LUT4 lut_inst_2264 (
  .F(lut_f_2264),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2264.INIT = 16'h8000;
LUT4 lut_inst_2265 (
  .F(lut_f_2265),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2265.INIT = 16'h8000;
LUT4 lut_inst_2266 (
  .F(lut_f_2266),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2266.INIT = 16'h8000;
LUT4 lut_inst_2267 (
  .F(lut_f_2267),
  .I0(lut_f_2264),
  .I1(lut_f_2265),
  .I2(lut_f_2266),
  .I3(gw_vcc)
);
defparam lut_inst_2267.INIT = 16'h8000;
LUT4 lut_inst_2268 (
  .F(lut_f_2268),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2268.INIT = 16'h8000;
LUT4 lut_inst_2269 (
  .F(lut_f_2269),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2269.INIT = 16'h8000;
LUT4 lut_inst_2270 (
  .F(lut_f_2270),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2270.INIT = 16'h8000;
LUT4 lut_inst_2271 (
  .F(lut_f_2271),
  .I0(lut_f_2268),
  .I1(lut_f_2269),
  .I2(lut_f_2270),
  .I3(gw_vcc)
);
defparam lut_inst_2271.INIT = 16'h8000;
LUT4 lut_inst_2272 (
  .F(lut_f_2272),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2272.INIT = 16'h8000;
LUT4 lut_inst_2273 (
  .F(lut_f_2273),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2273.INIT = 16'h8000;
LUT4 lut_inst_2274 (
  .F(lut_f_2274),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2274.INIT = 16'h8000;
LUT4 lut_inst_2275 (
  .F(lut_f_2275),
  .I0(lut_f_2272),
  .I1(lut_f_2273),
  .I2(lut_f_2274),
  .I3(gw_vcc)
);
defparam lut_inst_2275.INIT = 16'h8000;
LUT4 lut_inst_2276 (
  .F(lut_f_2276),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2276.INIT = 16'h8000;
LUT4 lut_inst_2277 (
  .F(lut_f_2277),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2277.INIT = 16'h8000;
LUT4 lut_inst_2278 (
  .F(lut_f_2278),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2278.INIT = 16'h8000;
LUT4 lut_inst_2279 (
  .F(lut_f_2279),
  .I0(lut_f_2276),
  .I1(lut_f_2277),
  .I2(lut_f_2278),
  .I3(gw_vcc)
);
defparam lut_inst_2279.INIT = 16'h8000;
LUT4 lut_inst_2280 (
  .F(lut_f_2280),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2280.INIT = 16'h8000;
LUT4 lut_inst_2281 (
  .F(lut_f_2281),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2281.INIT = 16'h8000;
LUT4 lut_inst_2282 (
  .F(lut_f_2282),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2282.INIT = 16'h8000;
LUT4 lut_inst_2283 (
  .F(lut_f_2283),
  .I0(lut_f_2280),
  .I1(lut_f_2281),
  .I2(lut_f_2282),
  .I3(gw_vcc)
);
defparam lut_inst_2283.INIT = 16'h8000;
LUT4 lut_inst_2284 (
  .F(lut_f_2284),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2284.INIT = 16'h8000;
LUT4 lut_inst_2285 (
  .F(lut_f_2285),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2285.INIT = 16'h8000;
LUT4 lut_inst_2286 (
  .F(lut_f_2286),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2286.INIT = 16'h8000;
LUT4 lut_inst_2287 (
  .F(lut_f_2287),
  .I0(lut_f_2284),
  .I1(lut_f_2285),
  .I2(lut_f_2286),
  .I3(gw_vcc)
);
defparam lut_inst_2287.INIT = 16'h8000;
LUT4 lut_inst_2288 (
  .F(lut_f_2288),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2288.INIT = 16'h8000;
LUT4 lut_inst_2289 (
  .F(lut_f_2289),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2289.INIT = 16'h8000;
LUT4 lut_inst_2290 (
  .F(lut_f_2290),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2290.INIT = 16'h8000;
LUT4 lut_inst_2291 (
  .F(lut_f_2291),
  .I0(lut_f_2288),
  .I1(lut_f_2289),
  .I2(lut_f_2290),
  .I3(gw_vcc)
);
defparam lut_inst_2291.INIT = 16'h8000;
LUT4 lut_inst_2292 (
  .F(lut_f_2292),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2292.INIT = 16'h8000;
LUT4 lut_inst_2293 (
  .F(lut_f_2293),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2293.INIT = 16'h8000;
LUT4 lut_inst_2294 (
  .F(lut_f_2294),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2294.INIT = 16'h8000;
LUT4 lut_inst_2295 (
  .F(lut_f_2295),
  .I0(lut_f_2292),
  .I1(lut_f_2293),
  .I2(lut_f_2294),
  .I3(gw_vcc)
);
defparam lut_inst_2295.INIT = 16'h8000;
LUT4 lut_inst_2296 (
  .F(lut_f_2296),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2296.INIT = 16'h8000;
LUT4 lut_inst_2297 (
  .F(lut_f_2297),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2297.INIT = 16'h8000;
LUT4 lut_inst_2298 (
  .F(lut_f_2298),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2298.INIT = 16'h8000;
LUT4 lut_inst_2299 (
  .F(lut_f_2299),
  .I0(lut_f_2296),
  .I1(lut_f_2297),
  .I2(lut_f_2298),
  .I3(gw_vcc)
);
defparam lut_inst_2299.INIT = 16'h8000;
LUT4 lut_inst_2300 (
  .F(lut_f_2300),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2300.INIT = 16'h8000;
LUT4 lut_inst_2301 (
  .F(lut_f_2301),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2301.INIT = 16'h8000;
LUT4 lut_inst_2302 (
  .F(lut_f_2302),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2302.INIT = 16'h8000;
LUT4 lut_inst_2303 (
  .F(lut_f_2303),
  .I0(lut_f_2300),
  .I1(lut_f_2301),
  .I2(lut_f_2302),
  .I3(gw_vcc)
);
defparam lut_inst_2303.INIT = 16'h8000;
LUT4 lut_inst_2304 (
  .F(lut_f_2304),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2304.INIT = 16'h8000;
LUT4 lut_inst_2305 (
  .F(lut_f_2305),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2305.INIT = 16'h8000;
LUT4 lut_inst_2306 (
  .F(lut_f_2306),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2306.INIT = 16'h8000;
LUT4 lut_inst_2307 (
  .F(lut_f_2307),
  .I0(lut_f_2304),
  .I1(lut_f_2305),
  .I2(lut_f_2306),
  .I3(gw_vcc)
);
defparam lut_inst_2307.INIT = 16'h8000;
LUT4 lut_inst_2308 (
  .F(lut_f_2308),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2308.INIT = 16'h8000;
LUT4 lut_inst_2309 (
  .F(lut_f_2309),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2309.INIT = 16'h8000;
LUT4 lut_inst_2310 (
  .F(lut_f_2310),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2310.INIT = 16'h8000;
LUT4 lut_inst_2311 (
  .F(lut_f_2311),
  .I0(lut_f_2308),
  .I1(lut_f_2309),
  .I2(lut_f_2310),
  .I3(gw_vcc)
);
defparam lut_inst_2311.INIT = 16'h8000;
LUT4 lut_inst_2312 (
  .F(lut_f_2312),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2312.INIT = 16'h8000;
LUT4 lut_inst_2313 (
  .F(lut_f_2313),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2313.INIT = 16'h8000;
LUT4 lut_inst_2314 (
  .F(lut_f_2314),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2314.INIT = 16'h8000;
LUT4 lut_inst_2315 (
  .F(lut_f_2315),
  .I0(lut_f_2312),
  .I1(lut_f_2313),
  .I2(lut_f_2314),
  .I3(gw_vcc)
);
defparam lut_inst_2315.INIT = 16'h8000;
LUT4 lut_inst_2316 (
  .F(lut_f_2316),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2316.INIT = 16'h8000;
LUT4 lut_inst_2317 (
  .F(lut_f_2317),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2317.INIT = 16'h8000;
LUT4 lut_inst_2318 (
  .F(lut_f_2318),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2318.INIT = 16'h8000;
LUT4 lut_inst_2319 (
  .F(lut_f_2319),
  .I0(lut_f_2316),
  .I1(lut_f_2317),
  .I2(lut_f_2318),
  .I3(gw_vcc)
);
defparam lut_inst_2319.INIT = 16'h8000;
LUT4 lut_inst_2320 (
  .F(lut_f_2320),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2320.INIT = 16'h8000;
LUT4 lut_inst_2321 (
  .F(lut_f_2321),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2321.INIT = 16'h8000;
LUT4 lut_inst_2322 (
  .F(lut_f_2322),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2322.INIT = 16'h8000;
LUT4 lut_inst_2323 (
  .F(lut_f_2323),
  .I0(lut_f_2320),
  .I1(lut_f_2321),
  .I2(lut_f_2322),
  .I3(gw_vcc)
);
defparam lut_inst_2323.INIT = 16'h8000;
LUT4 lut_inst_2324 (
  .F(lut_f_2324),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2324.INIT = 16'h8000;
LUT4 lut_inst_2325 (
  .F(lut_f_2325),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2325.INIT = 16'h8000;
LUT4 lut_inst_2326 (
  .F(lut_f_2326),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2326.INIT = 16'h8000;
LUT4 lut_inst_2327 (
  .F(lut_f_2327),
  .I0(lut_f_2324),
  .I1(lut_f_2325),
  .I2(lut_f_2326),
  .I3(gw_vcc)
);
defparam lut_inst_2327.INIT = 16'h8000;
LUT4 lut_inst_2328 (
  .F(lut_f_2328),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2328.INIT = 16'h8000;
LUT4 lut_inst_2329 (
  .F(lut_f_2329),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2329.INIT = 16'h8000;
LUT4 lut_inst_2330 (
  .F(lut_f_2330),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2330.INIT = 16'h8000;
LUT4 lut_inst_2331 (
  .F(lut_f_2331),
  .I0(lut_f_2328),
  .I1(lut_f_2329),
  .I2(lut_f_2330),
  .I3(gw_vcc)
);
defparam lut_inst_2331.INIT = 16'h8000;
LUT4 lut_inst_2332 (
  .F(lut_f_2332),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2332.INIT = 16'h8000;
LUT4 lut_inst_2333 (
  .F(lut_f_2333),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2333.INIT = 16'h8000;
LUT4 lut_inst_2334 (
  .F(lut_f_2334),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2334.INIT = 16'h8000;
LUT4 lut_inst_2335 (
  .F(lut_f_2335),
  .I0(lut_f_2332),
  .I1(lut_f_2333),
  .I2(lut_f_2334),
  .I3(gw_vcc)
);
defparam lut_inst_2335.INIT = 16'h8000;
LUT4 lut_inst_2336 (
  .F(lut_f_2336),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2336.INIT = 16'h8000;
LUT4 lut_inst_2337 (
  .F(lut_f_2337),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2337.INIT = 16'h8000;
LUT4 lut_inst_2338 (
  .F(lut_f_2338),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2338.INIT = 16'h8000;
LUT4 lut_inst_2339 (
  .F(lut_f_2339),
  .I0(lut_f_2336),
  .I1(lut_f_2337),
  .I2(lut_f_2338),
  .I3(gw_vcc)
);
defparam lut_inst_2339.INIT = 16'h8000;
LUT4 lut_inst_2340 (
  .F(lut_f_2340),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2340.INIT = 16'h8000;
LUT4 lut_inst_2341 (
  .F(lut_f_2341),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2341.INIT = 16'h8000;
LUT4 lut_inst_2342 (
  .F(lut_f_2342),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2342.INIT = 16'h8000;
LUT4 lut_inst_2343 (
  .F(lut_f_2343),
  .I0(lut_f_2340),
  .I1(lut_f_2341),
  .I2(lut_f_2342),
  .I3(gw_vcc)
);
defparam lut_inst_2343.INIT = 16'h8000;
LUT4 lut_inst_2344 (
  .F(lut_f_2344),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2344.INIT = 16'h8000;
LUT4 lut_inst_2345 (
  .F(lut_f_2345),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2345.INIT = 16'h8000;
LUT4 lut_inst_2346 (
  .F(lut_f_2346),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2346.INIT = 16'h8000;
LUT4 lut_inst_2347 (
  .F(lut_f_2347),
  .I0(lut_f_2344),
  .I1(lut_f_2345),
  .I2(lut_f_2346),
  .I3(gw_vcc)
);
defparam lut_inst_2347.INIT = 16'h8000;
LUT4 lut_inst_2348 (
  .F(lut_f_2348),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2348.INIT = 16'h8000;
LUT4 lut_inst_2349 (
  .F(lut_f_2349),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2349.INIT = 16'h8000;
LUT4 lut_inst_2350 (
  .F(lut_f_2350),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2350.INIT = 16'h8000;
LUT4 lut_inst_2351 (
  .F(lut_f_2351),
  .I0(lut_f_2348),
  .I1(lut_f_2349),
  .I2(lut_f_2350),
  .I3(gw_vcc)
);
defparam lut_inst_2351.INIT = 16'h8000;
LUT4 lut_inst_2352 (
  .F(lut_f_2352),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2352.INIT = 16'h8000;
LUT4 lut_inst_2353 (
  .F(lut_f_2353),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2353.INIT = 16'h8000;
LUT4 lut_inst_2354 (
  .F(lut_f_2354),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2354.INIT = 16'h8000;
LUT4 lut_inst_2355 (
  .F(lut_f_2355),
  .I0(lut_f_2352),
  .I1(lut_f_2353),
  .I2(lut_f_2354),
  .I3(gw_vcc)
);
defparam lut_inst_2355.INIT = 16'h8000;
LUT4 lut_inst_2356 (
  .F(lut_f_2356),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2356.INIT = 16'h8000;
LUT4 lut_inst_2357 (
  .F(lut_f_2357),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2357.INIT = 16'h8000;
LUT4 lut_inst_2358 (
  .F(lut_f_2358),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2358.INIT = 16'h8000;
LUT4 lut_inst_2359 (
  .F(lut_f_2359),
  .I0(lut_f_2356),
  .I1(lut_f_2357),
  .I2(lut_f_2358),
  .I3(gw_vcc)
);
defparam lut_inst_2359.INIT = 16'h8000;
LUT4 lut_inst_2360 (
  .F(lut_f_2360),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2360.INIT = 16'h8000;
LUT4 lut_inst_2361 (
  .F(lut_f_2361),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2361.INIT = 16'h8000;
LUT4 lut_inst_2362 (
  .F(lut_f_2362),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2362.INIT = 16'h8000;
LUT4 lut_inst_2363 (
  .F(lut_f_2363),
  .I0(lut_f_2360),
  .I1(lut_f_2361),
  .I2(lut_f_2362),
  .I3(gw_vcc)
);
defparam lut_inst_2363.INIT = 16'h8000;
LUT4 lut_inst_2364 (
  .F(lut_f_2364),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2364.INIT = 16'h8000;
LUT4 lut_inst_2365 (
  .F(lut_f_2365),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2365.INIT = 16'h8000;
LUT4 lut_inst_2366 (
  .F(lut_f_2366),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2366.INIT = 16'h8000;
LUT4 lut_inst_2367 (
  .F(lut_f_2367),
  .I0(lut_f_2364),
  .I1(lut_f_2365),
  .I2(lut_f_2366),
  .I3(gw_vcc)
);
defparam lut_inst_2367.INIT = 16'h8000;
LUT4 lut_inst_2368 (
  .F(lut_f_2368),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2368.INIT = 16'h8000;
LUT4 lut_inst_2369 (
  .F(lut_f_2369),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2369.INIT = 16'h8000;
LUT4 lut_inst_2370 (
  .F(lut_f_2370),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2370.INIT = 16'h8000;
LUT4 lut_inst_2371 (
  .F(lut_f_2371),
  .I0(lut_f_2368),
  .I1(lut_f_2369),
  .I2(lut_f_2370),
  .I3(gw_vcc)
);
defparam lut_inst_2371.INIT = 16'h8000;
LUT4 lut_inst_2372 (
  .F(lut_f_2372),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2372.INIT = 16'h8000;
LUT4 lut_inst_2373 (
  .F(lut_f_2373),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2373.INIT = 16'h8000;
LUT4 lut_inst_2374 (
  .F(lut_f_2374),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2374.INIT = 16'h8000;
LUT4 lut_inst_2375 (
  .F(lut_f_2375),
  .I0(lut_f_2372),
  .I1(lut_f_2373),
  .I2(lut_f_2374),
  .I3(gw_vcc)
);
defparam lut_inst_2375.INIT = 16'h8000;
LUT4 lut_inst_2376 (
  .F(lut_f_2376),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2376.INIT = 16'h8000;
LUT4 lut_inst_2377 (
  .F(lut_f_2377),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2377.INIT = 16'h8000;
LUT4 lut_inst_2378 (
  .F(lut_f_2378),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2378.INIT = 16'h8000;
LUT4 lut_inst_2379 (
  .F(lut_f_2379),
  .I0(lut_f_2376),
  .I1(lut_f_2377),
  .I2(lut_f_2378),
  .I3(gw_vcc)
);
defparam lut_inst_2379.INIT = 16'h8000;
LUT4 lut_inst_2380 (
  .F(lut_f_2380),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2380.INIT = 16'h8000;
LUT4 lut_inst_2381 (
  .F(lut_f_2381),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2381.INIT = 16'h8000;
LUT4 lut_inst_2382 (
  .F(lut_f_2382),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2382.INIT = 16'h8000;
LUT4 lut_inst_2383 (
  .F(lut_f_2383),
  .I0(lut_f_2380),
  .I1(lut_f_2381),
  .I2(lut_f_2382),
  .I3(gw_vcc)
);
defparam lut_inst_2383.INIT = 16'h8000;
LUT4 lut_inst_2384 (
  .F(lut_f_2384),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2384.INIT = 16'h8000;
LUT4 lut_inst_2385 (
  .F(lut_f_2385),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2385.INIT = 16'h8000;
LUT4 lut_inst_2386 (
  .F(lut_f_2386),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2386.INIT = 16'h8000;
LUT4 lut_inst_2387 (
  .F(lut_f_2387),
  .I0(lut_f_2384),
  .I1(lut_f_2385),
  .I2(lut_f_2386),
  .I3(gw_vcc)
);
defparam lut_inst_2387.INIT = 16'h8000;
LUT4 lut_inst_2388 (
  .F(lut_f_2388),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2388.INIT = 16'h8000;
LUT4 lut_inst_2389 (
  .F(lut_f_2389),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2389.INIT = 16'h8000;
LUT4 lut_inst_2390 (
  .F(lut_f_2390),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2390.INIT = 16'h8000;
LUT4 lut_inst_2391 (
  .F(lut_f_2391),
  .I0(lut_f_2388),
  .I1(lut_f_2389),
  .I2(lut_f_2390),
  .I3(gw_vcc)
);
defparam lut_inst_2391.INIT = 16'h8000;
LUT4 lut_inst_2392 (
  .F(lut_f_2392),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2392.INIT = 16'h8000;
LUT4 lut_inst_2393 (
  .F(lut_f_2393),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2393.INIT = 16'h8000;
LUT4 lut_inst_2394 (
  .F(lut_f_2394),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2394.INIT = 16'h8000;
LUT4 lut_inst_2395 (
  .F(lut_f_2395),
  .I0(lut_f_2392),
  .I1(lut_f_2393),
  .I2(lut_f_2394),
  .I3(gw_vcc)
);
defparam lut_inst_2395.INIT = 16'h8000;
LUT4 lut_inst_2396 (
  .F(lut_f_2396),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2396.INIT = 16'h8000;
LUT4 lut_inst_2397 (
  .F(lut_f_2397),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2397.INIT = 16'h8000;
LUT4 lut_inst_2398 (
  .F(lut_f_2398),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2398.INIT = 16'h8000;
LUT4 lut_inst_2399 (
  .F(lut_f_2399),
  .I0(lut_f_2396),
  .I1(lut_f_2397),
  .I2(lut_f_2398),
  .I3(gw_vcc)
);
defparam lut_inst_2399.INIT = 16'h8000;
LUT4 lut_inst_2400 (
  .F(lut_f_2400),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2400.INIT = 16'h8000;
LUT4 lut_inst_2401 (
  .F(lut_f_2401),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2401.INIT = 16'h8000;
LUT4 lut_inst_2402 (
  .F(lut_f_2402),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2402.INIT = 16'h8000;
LUT4 lut_inst_2403 (
  .F(lut_f_2403),
  .I0(lut_f_2400),
  .I1(lut_f_2401),
  .I2(lut_f_2402),
  .I3(gw_vcc)
);
defparam lut_inst_2403.INIT = 16'h8000;
LUT4 lut_inst_2404 (
  .F(lut_f_2404),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2404.INIT = 16'h8000;
LUT4 lut_inst_2405 (
  .F(lut_f_2405),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2405.INIT = 16'h8000;
LUT4 lut_inst_2406 (
  .F(lut_f_2406),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2406.INIT = 16'h8000;
LUT4 lut_inst_2407 (
  .F(lut_f_2407),
  .I0(lut_f_2404),
  .I1(lut_f_2405),
  .I2(lut_f_2406),
  .I3(gw_vcc)
);
defparam lut_inst_2407.INIT = 16'h8000;
LUT4 lut_inst_2408 (
  .F(lut_f_2408),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2408.INIT = 16'h8000;
LUT4 lut_inst_2409 (
  .F(lut_f_2409),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2409.INIT = 16'h8000;
LUT4 lut_inst_2410 (
  .F(lut_f_2410),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2410.INIT = 16'h8000;
LUT4 lut_inst_2411 (
  .F(lut_f_2411),
  .I0(lut_f_2408),
  .I1(lut_f_2409),
  .I2(lut_f_2410),
  .I3(gw_vcc)
);
defparam lut_inst_2411.INIT = 16'h8000;
LUT4 lut_inst_2412 (
  .F(lut_f_2412),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2412.INIT = 16'h8000;
LUT4 lut_inst_2413 (
  .F(lut_f_2413),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2413.INIT = 16'h8000;
LUT4 lut_inst_2414 (
  .F(lut_f_2414),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2414.INIT = 16'h8000;
LUT4 lut_inst_2415 (
  .F(lut_f_2415),
  .I0(lut_f_2412),
  .I1(lut_f_2413),
  .I2(lut_f_2414),
  .I3(gw_vcc)
);
defparam lut_inst_2415.INIT = 16'h8000;
LUT4 lut_inst_2416 (
  .F(lut_f_2416),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2416.INIT = 16'h8000;
LUT4 lut_inst_2417 (
  .F(lut_f_2417),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2417.INIT = 16'h8000;
LUT4 lut_inst_2418 (
  .F(lut_f_2418),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2418.INIT = 16'h8000;
LUT4 lut_inst_2419 (
  .F(lut_f_2419),
  .I0(lut_f_2416),
  .I1(lut_f_2417),
  .I2(lut_f_2418),
  .I3(gw_vcc)
);
defparam lut_inst_2419.INIT = 16'h8000;
LUT4 lut_inst_2420 (
  .F(lut_f_2420),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2420.INIT = 16'h8000;
LUT4 lut_inst_2421 (
  .F(lut_f_2421),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2421.INIT = 16'h8000;
LUT4 lut_inst_2422 (
  .F(lut_f_2422),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2422.INIT = 16'h8000;
LUT4 lut_inst_2423 (
  .F(lut_f_2423),
  .I0(lut_f_2420),
  .I1(lut_f_2421),
  .I2(lut_f_2422),
  .I3(gw_vcc)
);
defparam lut_inst_2423.INIT = 16'h8000;
LUT4 lut_inst_2424 (
  .F(lut_f_2424),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2424.INIT = 16'h8000;
LUT4 lut_inst_2425 (
  .F(lut_f_2425),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2425.INIT = 16'h8000;
LUT4 lut_inst_2426 (
  .F(lut_f_2426),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2426.INIT = 16'h8000;
LUT4 lut_inst_2427 (
  .F(lut_f_2427),
  .I0(lut_f_2424),
  .I1(lut_f_2425),
  .I2(lut_f_2426),
  .I3(gw_vcc)
);
defparam lut_inst_2427.INIT = 16'h8000;
LUT4 lut_inst_2428 (
  .F(lut_f_2428),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2428.INIT = 16'h8000;
LUT4 lut_inst_2429 (
  .F(lut_f_2429),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2429.INIT = 16'h8000;
LUT4 lut_inst_2430 (
  .F(lut_f_2430),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2430.INIT = 16'h8000;
LUT4 lut_inst_2431 (
  .F(lut_f_2431),
  .I0(lut_f_2428),
  .I1(lut_f_2429),
  .I2(lut_f_2430),
  .I3(gw_vcc)
);
defparam lut_inst_2431.INIT = 16'h8000;
LUT4 lut_inst_2432 (
  .F(lut_f_2432),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2432.INIT = 16'h8000;
LUT4 lut_inst_2433 (
  .F(lut_f_2433),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2433.INIT = 16'h8000;
LUT4 lut_inst_2434 (
  .F(lut_f_2434),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2434.INIT = 16'h8000;
LUT4 lut_inst_2435 (
  .F(lut_f_2435),
  .I0(lut_f_2432),
  .I1(lut_f_2433),
  .I2(lut_f_2434),
  .I3(gw_vcc)
);
defparam lut_inst_2435.INIT = 16'h8000;
LUT4 lut_inst_2436 (
  .F(lut_f_2436),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2436.INIT = 16'h8000;
LUT4 lut_inst_2437 (
  .F(lut_f_2437),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2437.INIT = 16'h8000;
LUT4 lut_inst_2438 (
  .F(lut_f_2438),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2438.INIT = 16'h8000;
LUT4 lut_inst_2439 (
  .F(lut_f_2439),
  .I0(lut_f_2436),
  .I1(lut_f_2437),
  .I2(lut_f_2438),
  .I3(gw_vcc)
);
defparam lut_inst_2439.INIT = 16'h8000;
LUT4 lut_inst_2440 (
  .F(lut_f_2440),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2440.INIT = 16'h8000;
LUT4 lut_inst_2441 (
  .F(lut_f_2441),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2441.INIT = 16'h8000;
LUT4 lut_inst_2442 (
  .F(lut_f_2442),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2442.INIT = 16'h8000;
LUT4 lut_inst_2443 (
  .F(lut_f_2443),
  .I0(lut_f_2440),
  .I1(lut_f_2441),
  .I2(lut_f_2442),
  .I3(gw_vcc)
);
defparam lut_inst_2443.INIT = 16'h8000;
LUT4 lut_inst_2444 (
  .F(lut_f_2444),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2444.INIT = 16'h8000;
LUT4 lut_inst_2445 (
  .F(lut_f_2445),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2445.INIT = 16'h8000;
LUT4 lut_inst_2446 (
  .F(lut_f_2446),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2446.INIT = 16'h8000;
LUT4 lut_inst_2447 (
  .F(lut_f_2447),
  .I0(lut_f_2444),
  .I1(lut_f_2445),
  .I2(lut_f_2446),
  .I3(gw_vcc)
);
defparam lut_inst_2447.INIT = 16'h8000;
LUT4 lut_inst_2448 (
  .F(lut_f_2448),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2448.INIT = 16'h8000;
LUT4 lut_inst_2449 (
  .F(lut_f_2449),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2449.INIT = 16'h8000;
LUT4 lut_inst_2450 (
  .F(lut_f_2450),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2450.INIT = 16'h8000;
LUT4 lut_inst_2451 (
  .F(lut_f_2451),
  .I0(lut_f_2448),
  .I1(lut_f_2449),
  .I2(lut_f_2450),
  .I3(gw_vcc)
);
defparam lut_inst_2451.INIT = 16'h8000;
LUT4 lut_inst_2452 (
  .F(lut_f_2452),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2452.INIT = 16'h8000;
LUT4 lut_inst_2453 (
  .F(lut_f_2453),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2453.INIT = 16'h8000;
LUT4 lut_inst_2454 (
  .F(lut_f_2454),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2454.INIT = 16'h8000;
LUT4 lut_inst_2455 (
  .F(lut_f_2455),
  .I0(lut_f_2452),
  .I1(lut_f_2453),
  .I2(lut_f_2454),
  .I3(gw_vcc)
);
defparam lut_inst_2455.INIT = 16'h8000;
LUT4 lut_inst_2456 (
  .F(lut_f_2456),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2456.INIT = 16'h8000;
LUT4 lut_inst_2457 (
  .F(lut_f_2457),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2457.INIT = 16'h8000;
LUT4 lut_inst_2458 (
  .F(lut_f_2458),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2458.INIT = 16'h8000;
LUT4 lut_inst_2459 (
  .F(lut_f_2459),
  .I0(lut_f_2456),
  .I1(lut_f_2457),
  .I2(lut_f_2458),
  .I3(gw_vcc)
);
defparam lut_inst_2459.INIT = 16'h8000;
LUT4 lut_inst_2460 (
  .F(lut_f_2460),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2460.INIT = 16'h8000;
LUT4 lut_inst_2461 (
  .F(lut_f_2461),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2461.INIT = 16'h8000;
LUT4 lut_inst_2462 (
  .F(lut_f_2462),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2462.INIT = 16'h8000;
LUT4 lut_inst_2463 (
  .F(lut_f_2463),
  .I0(lut_f_2460),
  .I1(lut_f_2461),
  .I2(lut_f_2462),
  .I3(gw_vcc)
);
defparam lut_inst_2463.INIT = 16'h8000;
LUT4 lut_inst_2464 (
  .F(lut_f_2464),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2464.INIT = 16'h8000;
LUT4 lut_inst_2465 (
  .F(lut_f_2465),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2465.INIT = 16'h8000;
LUT4 lut_inst_2466 (
  .F(lut_f_2466),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2466.INIT = 16'h8000;
LUT4 lut_inst_2467 (
  .F(lut_f_2467),
  .I0(lut_f_2464),
  .I1(lut_f_2465),
  .I2(lut_f_2466),
  .I3(gw_vcc)
);
defparam lut_inst_2467.INIT = 16'h8000;
LUT4 lut_inst_2468 (
  .F(lut_f_2468),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2468.INIT = 16'h8000;
LUT4 lut_inst_2469 (
  .F(lut_f_2469),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2469.INIT = 16'h8000;
LUT4 lut_inst_2470 (
  .F(lut_f_2470),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2470.INIT = 16'h8000;
LUT4 lut_inst_2471 (
  .F(lut_f_2471),
  .I0(lut_f_2468),
  .I1(lut_f_2469),
  .I2(lut_f_2470),
  .I3(gw_vcc)
);
defparam lut_inst_2471.INIT = 16'h8000;
LUT4 lut_inst_2472 (
  .F(lut_f_2472),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2472.INIT = 16'h8000;
LUT4 lut_inst_2473 (
  .F(lut_f_2473),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2473.INIT = 16'h8000;
LUT4 lut_inst_2474 (
  .F(lut_f_2474),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2474.INIT = 16'h8000;
LUT4 lut_inst_2475 (
  .F(lut_f_2475),
  .I0(lut_f_2472),
  .I1(lut_f_2473),
  .I2(lut_f_2474),
  .I3(gw_vcc)
);
defparam lut_inst_2475.INIT = 16'h8000;
LUT4 lut_inst_2476 (
  .F(lut_f_2476),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2476.INIT = 16'h8000;
LUT4 lut_inst_2477 (
  .F(lut_f_2477),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2477.INIT = 16'h8000;
LUT4 lut_inst_2478 (
  .F(lut_f_2478),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2478.INIT = 16'h8000;
LUT4 lut_inst_2479 (
  .F(lut_f_2479),
  .I0(lut_f_2476),
  .I1(lut_f_2477),
  .I2(lut_f_2478),
  .I3(gw_vcc)
);
defparam lut_inst_2479.INIT = 16'h8000;
LUT4 lut_inst_2480 (
  .F(lut_f_2480),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2480.INIT = 16'h8000;
LUT4 lut_inst_2481 (
  .F(lut_f_2481),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2481.INIT = 16'h8000;
LUT4 lut_inst_2482 (
  .F(lut_f_2482),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2482.INIT = 16'h8000;
LUT4 lut_inst_2483 (
  .F(lut_f_2483),
  .I0(lut_f_2480),
  .I1(lut_f_2481),
  .I2(lut_f_2482),
  .I3(gw_vcc)
);
defparam lut_inst_2483.INIT = 16'h8000;
LUT4 lut_inst_2484 (
  .F(lut_f_2484),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2484.INIT = 16'h8000;
LUT4 lut_inst_2485 (
  .F(lut_f_2485),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2485.INIT = 16'h8000;
LUT4 lut_inst_2486 (
  .F(lut_f_2486),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2486.INIT = 16'h8000;
LUT4 lut_inst_2487 (
  .F(lut_f_2487),
  .I0(lut_f_2484),
  .I1(lut_f_2485),
  .I2(lut_f_2486),
  .I3(gw_vcc)
);
defparam lut_inst_2487.INIT = 16'h8000;
LUT4 lut_inst_2488 (
  .F(lut_f_2488),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2488.INIT = 16'h8000;
LUT4 lut_inst_2489 (
  .F(lut_f_2489),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2489.INIT = 16'h8000;
LUT4 lut_inst_2490 (
  .F(lut_f_2490),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2490.INIT = 16'h8000;
LUT4 lut_inst_2491 (
  .F(lut_f_2491),
  .I0(lut_f_2488),
  .I1(lut_f_2489),
  .I2(lut_f_2490),
  .I3(gw_vcc)
);
defparam lut_inst_2491.INIT = 16'h8000;
LUT4 lut_inst_2492 (
  .F(lut_f_2492),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2492.INIT = 16'h8000;
LUT4 lut_inst_2493 (
  .F(lut_f_2493),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2493.INIT = 16'h8000;
LUT4 lut_inst_2494 (
  .F(lut_f_2494),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2494.INIT = 16'h8000;
LUT4 lut_inst_2495 (
  .F(lut_f_2495),
  .I0(lut_f_2492),
  .I1(lut_f_2493),
  .I2(lut_f_2494),
  .I3(gw_vcc)
);
defparam lut_inst_2495.INIT = 16'h8000;
LUT4 lut_inst_2496 (
  .F(lut_f_2496),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2496.INIT = 16'h8000;
LUT4 lut_inst_2497 (
  .F(lut_f_2497),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2497.INIT = 16'h8000;
LUT4 lut_inst_2498 (
  .F(lut_f_2498),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2498.INIT = 16'h8000;
LUT4 lut_inst_2499 (
  .F(lut_f_2499),
  .I0(lut_f_2496),
  .I1(lut_f_2497),
  .I2(lut_f_2498),
  .I3(gw_vcc)
);
defparam lut_inst_2499.INIT = 16'h8000;
LUT4 lut_inst_2500 (
  .F(lut_f_2500),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2500.INIT = 16'h8000;
LUT4 lut_inst_2501 (
  .F(lut_f_2501),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2501.INIT = 16'h8000;
LUT4 lut_inst_2502 (
  .F(lut_f_2502),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2502.INIT = 16'h8000;
LUT4 lut_inst_2503 (
  .F(lut_f_2503),
  .I0(lut_f_2500),
  .I1(lut_f_2501),
  .I2(lut_f_2502),
  .I3(gw_vcc)
);
defparam lut_inst_2503.INIT = 16'h8000;
LUT4 lut_inst_2504 (
  .F(lut_f_2504),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2504.INIT = 16'h8000;
LUT4 lut_inst_2505 (
  .F(lut_f_2505),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2505.INIT = 16'h8000;
LUT4 lut_inst_2506 (
  .F(lut_f_2506),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2506.INIT = 16'h8000;
LUT4 lut_inst_2507 (
  .F(lut_f_2507),
  .I0(lut_f_2504),
  .I1(lut_f_2505),
  .I2(lut_f_2506),
  .I3(gw_vcc)
);
defparam lut_inst_2507.INIT = 16'h8000;
LUT4 lut_inst_2508 (
  .F(lut_f_2508),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2508.INIT = 16'h8000;
LUT4 lut_inst_2509 (
  .F(lut_f_2509),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2509.INIT = 16'h8000;
LUT4 lut_inst_2510 (
  .F(lut_f_2510),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2510.INIT = 16'h8000;
LUT4 lut_inst_2511 (
  .F(lut_f_2511),
  .I0(lut_f_2508),
  .I1(lut_f_2509),
  .I2(lut_f_2510),
  .I3(gw_vcc)
);
defparam lut_inst_2511.INIT = 16'h8000;
LUT4 lut_inst_2512 (
  .F(lut_f_2512),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2512.INIT = 16'h8000;
LUT4 lut_inst_2513 (
  .F(lut_f_2513),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2513.INIT = 16'h8000;
LUT4 lut_inst_2514 (
  .F(lut_f_2514),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2514.INIT = 16'h8000;
LUT4 lut_inst_2515 (
  .F(lut_f_2515),
  .I0(lut_f_2512),
  .I1(lut_f_2513),
  .I2(lut_f_2514),
  .I3(gw_vcc)
);
defparam lut_inst_2515.INIT = 16'h8000;
LUT4 lut_inst_2516 (
  .F(lut_f_2516),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2516.INIT = 16'h8000;
LUT4 lut_inst_2517 (
  .F(lut_f_2517),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2517.INIT = 16'h8000;
LUT4 lut_inst_2518 (
  .F(lut_f_2518),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2518.INIT = 16'h8000;
LUT4 lut_inst_2519 (
  .F(lut_f_2519),
  .I0(lut_f_2516),
  .I1(lut_f_2517),
  .I2(lut_f_2518),
  .I3(gw_vcc)
);
defparam lut_inst_2519.INIT = 16'h8000;
LUT4 lut_inst_2520 (
  .F(lut_f_2520),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2520.INIT = 16'h8000;
LUT4 lut_inst_2521 (
  .F(lut_f_2521),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2521.INIT = 16'h8000;
LUT4 lut_inst_2522 (
  .F(lut_f_2522),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2522.INIT = 16'h8000;
LUT4 lut_inst_2523 (
  .F(lut_f_2523),
  .I0(lut_f_2520),
  .I1(lut_f_2521),
  .I2(lut_f_2522),
  .I3(gw_vcc)
);
defparam lut_inst_2523.INIT = 16'h8000;
LUT4 lut_inst_2524 (
  .F(lut_f_2524),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2524.INIT = 16'h8000;
LUT4 lut_inst_2525 (
  .F(lut_f_2525),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2525.INIT = 16'h8000;
LUT4 lut_inst_2526 (
  .F(lut_f_2526),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2526.INIT = 16'h8000;
LUT4 lut_inst_2527 (
  .F(lut_f_2527),
  .I0(lut_f_2524),
  .I1(lut_f_2525),
  .I2(lut_f_2526),
  .I3(gw_vcc)
);
defparam lut_inst_2527.INIT = 16'h8000;
LUT4 lut_inst_2528 (
  .F(lut_f_2528),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2528.INIT = 16'h8000;
LUT4 lut_inst_2529 (
  .F(lut_f_2529),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2529.INIT = 16'h8000;
LUT4 lut_inst_2530 (
  .F(lut_f_2530),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2530.INIT = 16'h8000;
LUT4 lut_inst_2531 (
  .F(lut_f_2531),
  .I0(lut_f_2528),
  .I1(lut_f_2529),
  .I2(lut_f_2530),
  .I3(gw_vcc)
);
defparam lut_inst_2531.INIT = 16'h8000;
LUT4 lut_inst_2532 (
  .F(lut_f_2532),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2532.INIT = 16'h8000;
LUT4 lut_inst_2533 (
  .F(lut_f_2533),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2533.INIT = 16'h8000;
LUT4 lut_inst_2534 (
  .F(lut_f_2534),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2534.INIT = 16'h8000;
LUT4 lut_inst_2535 (
  .F(lut_f_2535),
  .I0(lut_f_2532),
  .I1(lut_f_2533),
  .I2(lut_f_2534),
  .I3(gw_vcc)
);
defparam lut_inst_2535.INIT = 16'h8000;
LUT4 lut_inst_2536 (
  .F(lut_f_2536),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2536.INIT = 16'h8000;
LUT4 lut_inst_2537 (
  .F(lut_f_2537),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2537.INIT = 16'h8000;
LUT4 lut_inst_2538 (
  .F(lut_f_2538),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2538.INIT = 16'h8000;
LUT4 lut_inst_2539 (
  .F(lut_f_2539),
  .I0(lut_f_2536),
  .I1(lut_f_2537),
  .I2(lut_f_2538),
  .I3(gw_vcc)
);
defparam lut_inst_2539.INIT = 16'h8000;
LUT4 lut_inst_2540 (
  .F(lut_f_2540),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2540.INIT = 16'h8000;
LUT4 lut_inst_2541 (
  .F(lut_f_2541),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2541.INIT = 16'h8000;
LUT4 lut_inst_2542 (
  .F(lut_f_2542),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2542.INIT = 16'h8000;
LUT4 lut_inst_2543 (
  .F(lut_f_2543),
  .I0(lut_f_2540),
  .I1(lut_f_2541),
  .I2(lut_f_2542),
  .I3(gw_vcc)
);
defparam lut_inst_2543.INIT = 16'h8000;
LUT4 lut_inst_2544 (
  .F(lut_f_2544),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2544.INIT = 16'h8000;
LUT4 lut_inst_2545 (
  .F(lut_f_2545),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2545.INIT = 16'h8000;
LUT4 lut_inst_2546 (
  .F(lut_f_2546),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2546.INIT = 16'h8000;
LUT4 lut_inst_2547 (
  .F(lut_f_2547),
  .I0(lut_f_2544),
  .I1(lut_f_2545),
  .I2(lut_f_2546),
  .I3(gw_vcc)
);
defparam lut_inst_2547.INIT = 16'h8000;
LUT4 lut_inst_2548 (
  .F(lut_f_2548),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2548.INIT = 16'h8000;
LUT4 lut_inst_2549 (
  .F(lut_f_2549),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2549.INIT = 16'h8000;
LUT4 lut_inst_2550 (
  .F(lut_f_2550),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2550.INIT = 16'h8000;
LUT4 lut_inst_2551 (
  .F(lut_f_2551),
  .I0(lut_f_2548),
  .I1(lut_f_2549),
  .I2(lut_f_2550),
  .I3(gw_vcc)
);
defparam lut_inst_2551.INIT = 16'h8000;
LUT4 lut_inst_2552 (
  .F(lut_f_2552),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2552.INIT = 16'h8000;
LUT4 lut_inst_2553 (
  .F(lut_f_2553),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2553.INIT = 16'h8000;
LUT4 lut_inst_2554 (
  .F(lut_f_2554),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2554.INIT = 16'h8000;
LUT4 lut_inst_2555 (
  .F(lut_f_2555),
  .I0(lut_f_2552),
  .I1(lut_f_2553),
  .I2(lut_f_2554),
  .I3(gw_vcc)
);
defparam lut_inst_2555.INIT = 16'h8000;
LUT4 lut_inst_2556 (
  .F(lut_f_2556),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2556.INIT = 16'h8000;
LUT4 lut_inst_2557 (
  .F(lut_f_2557),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2557.INIT = 16'h8000;
LUT4 lut_inst_2558 (
  .F(lut_f_2558),
  .I0(ad11_inv),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2558.INIT = 16'h8000;
LUT4 lut_inst_2559 (
  .F(lut_f_2559),
  .I0(lut_f_2556),
  .I1(lut_f_2557),
  .I2(lut_f_2558),
  .I3(gw_vcc)
);
defparam lut_inst_2559.INIT = 16'h8000;
LUT4 lut_inst_2560 (
  .F(lut_f_2560),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2560.INIT = 16'h8000;
LUT4 lut_inst_2561 (
  .F(lut_f_2561),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2561.INIT = 16'h8000;
LUT4 lut_inst_2562 (
  .F(lut_f_2562),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2562.INIT = 16'h8000;
LUT4 lut_inst_2563 (
  .F(lut_f_2563),
  .I0(lut_f_2560),
  .I1(lut_f_2561),
  .I2(lut_f_2562),
  .I3(gw_vcc)
);
defparam lut_inst_2563.INIT = 16'h8000;
LUT4 lut_inst_2564 (
  .F(lut_f_2564),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2564.INIT = 16'h8000;
LUT4 lut_inst_2565 (
  .F(lut_f_2565),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2565.INIT = 16'h8000;
LUT4 lut_inst_2566 (
  .F(lut_f_2566),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2566.INIT = 16'h8000;
LUT4 lut_inst_2567 (
  .F(lut_f_2567),
  .I0(lut_f_2564),
  .I1(lut_f_2565),
  .I2(lut_f_2566),
  .I3(gw_vcc)
);
defparam lut_inst_2567.INIT = 16'h8000;
LUT4 lut_inst_2568 (
  .F(lut_f_2568),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2568.INIT = 16'h8000;
LUT4 lut_inst_2569 (
  .F(lut_f_2569),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2569.INIT = 16'h8000;
LUT4 lut_inst_2570 (
  .F(lut_f_2570),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2570.INIT = 16'h8000;
LUT4 lut_inst_2571 (
  .F(lut_f_2571),
  .I0(lut_f_2568),
  .I1(lut_f_2569),
  .I2(lut_f_2570),
  .I3(gw_vcc)
);
defparam lut_inst_2571.INIT = 16'h8000;
LUT4 lut_inst_2572 (
  .F(lut_f_2572),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2572.INIT = 16'h8000;
LUT4 lut_inst_2573 (
  .F(lut_f_2573),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2573.INIT = 16'h8000;
LUT4 lut_inst_2574 (
  .F(lut_f_2574),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2574.INIT = 16'h8000;
LUT4 lut_inst_2575 (
  .F(lut_f_2575),
  .I0(lut_f_2572),
  .I1(lut_f_2573),
  .I2(lut_f_2574),
  .I3(gw_vcc)
);
defparam lut_inst_2575.INIT = 16'h8000;
LUT4 lut_inst_2576 (
  .F(lut_f_2576),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2576.INIT = 16'h8000;
LUT4 lut_inst_2577 (
  .F(lut_f_2577),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2577.INIT = 16'h8000;
LUT4 lut_inst_2578 (
  .F(lut_f_2578),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2578.INIT = 16'h8000;
LUT4 lut_inst_2579 (
  .F(lut_f_2579),
  .I0(lut_f_2576),
  .I1(lut_f_2577),
  .I2(lut_f_2578),
  .I3(gw_vcc)
);
defparam lut_inst_2579.INIT = 16'h8000;
LUT4 lut_inst_2580 (
  .F(lut_f_2580),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2580.INIT = 16'h8000;
LUT4 lut_inst_2581 (
  .F(lut_f_2581),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2581.INIT = 16'h8000;
LUT4 lut_inst_2582 (
  .F(lut_f_2582),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2582.INIT = 16'h8000;
LUT4 lut_inst_2583 (
  .F(lut_f_2583),
  .I0(lut_f_2580),
  .I1(lut_f_2581),
  .I2(lut_f_2582),
  .I3(gw_vcc)
);
defparam lut_inst_2583.INIT = 16'h8000;
LUT4 lut_inst_2584 (
  .F(lut_f_2584),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2584.INIT = 16'h8000;
LUT4 lut_inst_2585 (
  .F(lut_f_2585),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2585.INIT = 16'h8000;
LUT4 lut_inst_2586 (
  .F(lut_f_2586),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2586.INIT = 16'h8000;
LUT4 lut_inst_2587 (
  .F(lut_f_2587),
  .I0(lut_f_2584),
  .I1(lut_f_2585),
  .I2(lut_f_2586),
  .I3(gw_vcc)
);
defparam lut_inst_2587.INIT = 16'h8000;
LUT4 lut_inst_2588 (
  .F(lut_f_2588),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2588.INIT = 16'h8000;
LUT4 lut_inst_2589 (
  .F(lut_f_2589),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2589.INIT = 16'h8000;
LUT4 lut_inst_2590 (
  .F(lut_f_2590),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2590.INIT = 16'h8000;
LUT4 lut_inst_2591 (
  .F(lut_f_2591),
  .I0(lut_f_2588),
  .I1(lut_f_2589),
  .I2(lut_f_2590),
  .I3(gw_vcc)
);
defparam lut_inst_2591.INIT = 16'h8000;
LUT4 lut_inst_2592 (
  .F(lut_f_2592),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2592.INIT = 16'h8000;
LUT4 lut_inst_2593 (
  .F(lut_f_2593),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2593.INIT = 16'h8000;
LUT4 lut_inst_2594 (
  .F(lut_f_2594),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2594.INIT = 16'h8000;
LUT4 lut_inst_2595 (
  .F(lut_f_2595),
  .I0(lut_f_2592),
  .I1(lut_f_2593),
  .I2(lut_f_2594),
  .I3(gw_vcc)
);
defparam lut_inst_2595.INIT = 16'h8000;
LUT4 lut_inst_2596 (
  .F(lut_f_2596),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2596.INIT = 16'h8000;
LUT4 lut_inst_2597 (
  .F(lut_f_2597),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2597.INIT = 16'h8000;
LUT4 lut_inst_2598 (
  .F(lut_f_2598),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2598.INIT = 16'h8000;
LUT4 lut_inst_2599 (
  .F(lut_f_2599),
  .I0(lut_f_2596),
  .I1(lut_f_2597),
  .I2(lut_f_2598),
  .I3(gw_vcc)
);
defparam lut_inst_2599.INIT = 16'h8000;
LUT4 lut_inst_2600 (
  .F(lut_f_2600),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2600.INIT = 16'h8000;
LUT4 lut_inst_2601 (
  .F(lut_f_2601),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2601.INIT = 16'h8000;
LUT4 lut_inst_2602 (
  .F(lut_f_2602),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2602.INIT = 16'h8000;
LUT4 lut_inst_2603 (
  .F(lut_f_2603),
  .I0(lut_f_2600),
  .I1(lut_f_2601),
  .I2(lut_f_2602),
  .I3(gw_vcc)
);
defparam lut_inst_2603.INIT = 16'h8000;
LUT4 lut_inst_2604 (
  .F(lut_f_2604),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2604.INIT = 16'h8000;
LUT4 lut_inst_2605 (
  .F(lut_f_2605),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2605.INIT = 16'h8000;
LUT4 lut_inst_2606 (
  .F(lut_f_2606),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2606.INIT = 16'h8000;
LUT4 lut_inst_2607 (
  .F(lut_f_2607),
  .I0(lut_f_2604),
  .I1(lut_f_2605),
  .I2(lut_f_2606),
  .I3(gw_vcc)
);
defparam lut_inst_2607.INIT = 16'h8000;
LUT4 lut_inst_2608 (
  .F(lut_f_2608),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2608.INIT = 16'h8000;
LUT4 lut_inst_2609 (
  .F(lut_f_2609),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2609.INIT = 16'h8000;
LUT4 lut_inst_2610 (
  .F(lut_f_2610),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2610.INIT = 16'h8000;
LUT4 lut_inst_2611 (
  .F(lut_f_2611),
  .I0(lut_f_2608),
  .I1(lut_f_2609),
  .I2(lut_f_2610),
  .I3(gw_vcc)
);
defparam lut_inst_2611.INIT = 16'h8000;
LUT4 lut_inst_2612 (
  .F(lut_f_2612),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2612.INIT = 16'h8000;
LUT4 lut_inst_2613 (
  .F(lut_f_2613),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2613.INIT = 16'h8000;
LUT4 lut_inst_2614 (
  .F(lut_f_2614),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2614.INIT = 16'h8000;
LUT4 lut_inst_2615 (
  .F(lut_f_2615),
  .I0(lut_f_2612),
  .I1(lut_f_2613),
  .I2(lut_f_2614),
  .I3(gw_vcc)
);
defparam lut_inst_2615.INIT = 16'h8000;
LUT4 lut_inst_2616 (
  .F(lut_f_2616),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2616.INIT = 16'h8000;
LUT4 lut_inst_2617 (
  .F(lut_f_2617),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2617.INIT = 16'h8000;
LUT4 lut_inst_2618 (
  .F(lut_f_2618),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2618.INIT = 16'h8000;
LUT4 lut_inst_2619 (
  .F(lut_f_2619),
  .I0(lut_f_2616),
  .I1(lut_f_2617),
  .I2(lut_f_2618),
  .I3(gw_vcc)
);
defparam lut_inst_2619.INIT = 16'h8000;
LUT4 lut_inst_2620 (
  .F(lut_f_2620),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2620.INIT = 16'h8000;
LUT4 lut_inst_2621 (
  .F(lut_f_2621),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2621.INIT = 16'h8000;
LUT4 lut_inst_2622 (
  .F(lut_f_2622),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2622.INIT = 16'h8000;
LUT4 lut_inst_2623 (
  .F(lut_f_2623),
  .I0(lut_f_2620),
  .I1(lut_f_2621),
  .I2(lut_f_2622),
  .I3(gw_vcc)
);
defparam lut_inst_2623.INIT = 16'h8000;
LUT4 lut_inst_2624 (
  .F(lut_f_2624),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2624.INIT = 16'h8000;
LUT4 lut_inst_2625 (
  .F(lut_f_2625),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2625.INIT = 16'h8000;
LUT4 lut_inst_2626 (
  .F(lut_f_2626),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2626.INIT = 16'h8000;
LUT4 lut_inst_2627 (
  .F(lut_f_2627),
  .I0(lut_f_2624),
  .I1(lut_f_2625),
  .I2(lut_f_2626),
  .I3(gw_vcc)
);
defparam lut_inst_2627.INIT = 16'h8000;
LUT4 lut_inst_2628 (
  .F(lut_f_2628),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2628.INIT = 16'h8000;
LUT4 lut_inst_2629 (
  .F(lut_f_2629),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2629.INIT = 16'h8000;
LUT4 lut_inst_2630 (
  .F(lut_f_2630),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2630.INIT = 16'h8000;
LUT4 lut_inst_2631 (
  .F(lut_f_2631),
  .I0(lut_f_2628),
  .I1(lut_f_2629),
  .I2(lut_f_2630),
  .I3(gw_vcc)
);
defparam lut_inst_2631.INIT = 16'h8000;
LUT4 lut_inst_2632 (
  .F(lut_f_2632),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2632.INIT = 16'h8000;
LUT4 lut_inst_2633 (
  .F(lut_f_2633),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2633.INIT = 16'h8000;
LUT4 lut_inst_2634 (
  .F(lut_f_2634),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2634.INIT = 16'h8000;
LUT4 lut_inst_2635 (
  .F(lut_f_2635),
  .I0(lut_f_2632),
  .I1(lut_f_2633),
  .I2(lut_f_2634),
  .I3(gw_vcc)
);
defparam lut_inst_2635.INIT = 16'h8000;
LUT4 lut_inst_2636 (
  .F(lut_f_2636),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2636.INIT = 16'h8000;
LUT4 lut_inst_2637 (
  .F(lut_f_2637),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2637.INIT = 16'h8000;
LUT4 lut_inst_2638 (
  .F(lut_f_2638),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2638.INIT = 16'h8000;
LUT4 lut_inst_2639 (
  .F(lut_f_2639),
  .I0(lut_f_2636),
  .I1(lut_f_2637),
  .I2(lut_f_2638),
  .I3(gw_vcc)
);
defparam lut_inst_2639.INIT = 16'h8000;
LUT4 lut_inst_2640 (
  .F(lut_f_2640),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2640.INIT = 16'h8000;
LUT4 lut_inst_2641 (
  .F(lut_f_2641),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2641.INIT = 16'h8000;
LUT4 lut_inst_2642 (
  .F(lut_f_2642),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2642.INIT = 16'h8000;
LUT4 lut_inst_2643 (
  .F(lut_f_2643),
  .I0(lut_f_2640),
  .I1(lut_f_2641),
  .I2(lut_f_2642),
  .I3(gw_vcc)
);
defparam lut_inst_2643.INIT = 16'h8000;
LUT4 lut_inst_2644 (
  .F(lut_f_2644),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2644.INIT = 16'h8000;
LUT4 lut_inst_2645 (
  .F(lut_f_2645),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2645.INIT = 16'h8000;
LUT4 lut_inst_2646 (
  .F(lut_f_2646),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2646.INIT = 16'h8000;
LUT4 lut_inst_2647 (
  .F(lut_f_2647),
  .I0(lut_f_2644),
  .I1(lut_f_2645),
  .I2(lut_f_2646),
  .I3(gw_vcc)
);
defparam lut_inst_2647.INIT = 16'h8000;
LUT4 lut_inst_2648 (
  .F(lut_f_2648),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2648.INIT = 16'h8000;
LUT4 lut_inst_2649 (
  .F(lut_f_2649),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2649.INIT = 16'h8000;
LUT4 lut_inst_2650 (
  .F(lut_f_2650),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2650.INIT = 16'h8000;
LUT4 lut_inst_2651 (
  .F(lut_f_2651),
  .I0(lut_f_2648),
  .I1(lut_f_2649),
  .I2(lut_f_2650),
  .I3(gw_vcc)
);
defparam lut_inst_2651.INIT = 16'h8000;
LUT4 lut_inst_2652 (
  .F(lut_f_2652),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2652.INIT = 16'h8000;
LUT4 lut_inst_2653 (
  .F(lut_f_2653),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2653.INIT = 16'h8000;
LUT4 lut_inst_2654 (
  .F(lut_f_2654),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2654.INIT = 16'h8000;
LUT4 lut_inst_2655 (
  .F(lut_f_2655),
  .I0(lut_f_2652),
  .I1(lut_f_2653),
  .I2(lut_f_2654),
  .I3(gw_vcc)
);
defparam lut_inst_2655.INIT = 16'h8000;
LUT4 lut_inst_2656 (
  .F(lut_f_2656),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2656.INIT = 16'h8000;
LUT4 lut_inst_2657 (
  .F(lut_f_2657),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2657.INIT = 16'h8000;
LUT4 lut_inst_2658 (
  .F(lut_f_2658),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2658.INIT = 16'h8000;
LUT4 lut_inst_2659 (
  .F(lut_f_2659),
  .I0(lut_f_2656),
  .I1(lut_f_2657),
  .I2(lut_f_2658),
  .I3(gw_vcc)
);
defparam lut_inst_2659.INIT = 16'h8000;
LUT4 lut_inst_2660 (
  .F(lut_f_2660),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2660.INIT = 16'h8000;
LUT4 lut_inst_2661 (
  .F(lut_f_2661),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2661.INIT = 16'h8000;
LUT4 lut_inst_2662 (
  .F(lut_f_2662),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2662.INIT = 16'h8000;
LUT4 lut_inst_2663 (
  .F(lut_f_2663),
  .I0(lut_f_2660),
  .I1(lut_f_2661),
  .I2(lut_f_2662),
  .I3(gw_vcc)
);
defparam lut_inst_2663.INIT = 16'h8000;
LUT4 lut_inst_2664 (
  .F(lut_f_2664),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2664.INIT = 16'h8000;
LUT4 lut_inst_2665 (
  .F(lut_f_2665),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2665.INIT = 16'h8000;
LUT4 lut_inst_2666 (
  .F(lut_f_2666),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2666.INIT = 16'h8000;
LUT4 lut_inst_2667 (
  .F(lut_f_2667),
  .I0(lut_f_2664),
  .I1(lut_f_2665),
  .I2(lut_f_2666),
  .I3(gw_vcc)
);
defparam lut_inst_2667.INIT = 16'h8000;
LUT4 lut_inst_2668 (
  .F(lut_f_2668),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2668.INIT = 16'h8000;
LUT4 lut_inst_2669 (
  .F(lut_f_2669),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2669.INIT = 16'h8000;
LUT4 lut_inst_2670 (
  .F(lut_f_2670),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2670.INIT = 16'h8000;
LUT4 lut_inst_2671 (
  .F(lut_f_2671),
  .I0(lut_f_2668),
  .I1(lut_f_2669),
  .I2(lut_f_2670),
  .I3(gw_vcc)
);
defparam lut_inst_2671.INIT = 16'h8000;
LUT4 lut_inst_2672 (
  .F(lut_f_2672),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2672.INIT = 16'h8000;
LUT4 lut_inst_2673 (
  .F(lut_f_2673),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2673.INIT = 16'h8000;
LUT4 lut_inst_2674 (
  .F(lut_f_2674),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2674.INIT = 16'h8000;
LUT4 lut_inst_2675 (
  .F(lut_f_2675),
  .I0(lut_f_2672),
  .I1(lut_f_2673),
  .I2(lut_f_2674),
  .I3(gw_vcc)
);
defparam lut_inst_2675.INIT = 16'h8000;
LUT4 lut_inst_2676 (
  .F(lut_f_2676),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2676.INIT = 16'h8000;
LUT4 lut_inst_2677 (
  .F(lut_f_2677),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2677.INIT = 16'h8000;
LUT4 lut_inst_2678 (
  .F(lut_f_2678),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2678.INIT = 16'h8000;
LUT4 lut_inst_2679 (
  .F(lut_f_2679),
  .I0(lut_f_2676),
  .I1(lut_f_2677),
  .I2(lut_f_2678),
  .I3(gw_vcc)
);
defparam lut_inst_2679.INIT = 16'h8000;
LUT4 lut_inst_2680 (
  .F(lut_f_2680),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2680.INIT = 16'h8000;
LUT4 lut_inst_2681 (
  .F(lut_f_2681),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2681.INIT = 16'h8000;
LUT4 lut_inst_2682 (
  .F(lut_f_2682),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2682.INIT = 16'h8000;
LUT4 lut_inst_2683 (
  .F(lut_f_2683),
  .I0(lut_f_2680),
  .I1(lut_f_2681),
  .I2(lut_f_2682),
  .I3(gw_vcc)
);
defparam lut_inst_2683.INIT = 16'h8000;
LUT4 lut_inst_2684 (
  .F(lut_f_2684),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2684.INIT = 16'h8000;
LUT4 lut_inst_2685 (
  .F(lut_f_2685),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_2685.INIT = 16'h8000;
LUT4 lut_inst_2686 (
  .F(lut_f_2686),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2686.INIT = 16'h8000;
LUT4 lut_inst_2687 (
  .F(lut_f_2687),
  .I0(lut_f_2684),
  .I1(lut_f_2685),
  .I2(lut_f_2686),
  .I3(gw_vcc)
);
defparam lut_inst_2687.INIT = 16'h8000;
LUT4 lut_inst_2688 (
  .F(lut_f_2688),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2688.INIT = 16'h8000;
LUT4 lut_inst_2689 (
  .F(lut_f_2689),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2689.INIT = 16'h8000;
LUT4 lut_inst_2690 (
  .F(lut_f_2690),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2690.INIT = 16'h8000;
LUT4 lut_inst_2691 (
  .F(lut_f_2691),
  .I0(lut_f_2688),
  .I1(lut_f_2689),
  .I2(lut_f_2690),
  .I3(gw_vcc)
);
defparam lut_inst_2691.INIT = 16'h8000;
LUT4 lut_inst_2692 (
  .F(lut_f_2692),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2692.INIT = 16'h8000;
LUT4 lut_inst_2693 (
  .F(lut_f_2693),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2693.INIT = 16'h8000;
LUT4 lut_inst_2694 (
  .F(lut_f_2694),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2694.INIT = 16'h8000;
LUT4 lut_inst_2695 (
  .F(lut_f_2695),
  .I0(lut_f_2692),
  .I1(lut_f_2693),
  .I2(lut_f_2694),
  .I3(gw_vcc)
);
defparam lut_inst_2695.INIT = 16'h8000;
LUT4 lut_inst_2696 (
  .F(lut_f_2696),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2696.INIT = 16'h8000;
LUT4 lut_inst_2697 (
  .F(lut_f_2697),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2697.INIT = 16'h8000;
LUT4 lut_inst_2698 (
  .F(lut_f_2698),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2698.INIT = 16'h8000;
LUT4 lut_inst_2699 (
  .F(lut_f_2699),
  .I0(lut_f_2696),
  .I1(lut_f_2697),
  .I2(lut_f_2698),
  .I3(gw_vcc)
);
defparam lut_inst_2699.INIT = 16'h8000;
LUT4 lut_inst_2700 (
  .F(lut_f_2700),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2700.INIT = 16'h8000;
LUT4 lut_inst_2701 (
  .F(lut_f_2701),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2701.INIT = 16'h8000;
LUT4 lut_inst_2702 (
  .F(lut_f_2702),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2702.INIT = 16'h8000;
LUT4 lut_inst_2703 (
  .F(lut_f_2703),
  .I0(lut_f_2700),
  .I1(lut_f_2701),
  .I2(lut_f_2702),
  .I3(gw_vcc)
);
defparam lut_inst_2703.INIT = 16'h8000;
LUT4 lut_inst_2704 (
  .F(lut_f_2704),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2704.INIT = 16'h8000;
LUT4 lut_inst_2705 (
  .F(lut_f_2705),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2705.INIT = 16'h8000;
LUT4 lut_inst_2706 (
  .F(lut_f_2706),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2706.INIT = 16'h8000;
LUT4 lut_inst_2707 (
  .F(lut_f_2707),
  .I0(lut_f_2704),
  .I1(lut_f_2705),
  .I2(lut_f_2706),
  .I3(gw_vcc)
);
defparam lut_inst_2707.INIT = 16'h8000;
LUT4 lut_inst_2708 (
  .F(lut_f_2708),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2708.INIT = 16'h8000;
LUT4 lut_inst_2709 (
  .F(lut_f_2709),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2709.INIT = 16'h8000;
LUT4 lut_inst_2710 (
  .F(lut_f_2710),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2710.INIT = 16'h8000;
LUT4 lut_inst_2711 (
  .F(lut_f_2711),
  .I0(lut_f_2708),
  .I1(lut_f_2709),
  .I2(lut_f_2710),
  .I3(gw_vcc)
);
defparam lut_inst_2711.INIT = 16'h8000;
LUT4 lut_inst_2712 (
  .F(lut_f_2712),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2712.INIT = 16'h8000;
LUT4 lut_inst_2713 (
  .F(lut_f_2713),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2713.INIT = 16'h8000;
LUT4 lut_inst_2714 (
  .F(lut_f_2714),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2714.INIT = 16'h8000;
LUT4 lut_inst_2715 (
  .F(lut_f_2715),
  .I0(lut_f_2712),
  .I1(lut_f_2713),
  .I2(lut_f_2714),
  .I3(gw_vcc)
);
defparam lut_inst_2715.INIT = 16'h8000;
LUT4 lut_inst_2716 (
  .F(lut_f_2716),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2716.INIT = 16'h8000;
LUT4 lut_inst_2717 (
  .F(lut_f_2717),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2717.INIT = 16'h8000;
LUT4 lut_inst_2718 (
  .F(lut_f_2718),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2718.INIT = 16'h8000;
LUT4 lut_inst_2719 (
  .F(lut_f_2719),
  .I0(lut_f_2716),
  .I1(lut_f_2717),
  .I2(lut_f_2718),
  .I3(gw_vcc)
);
defparam lut_inst_2719.INIT = 16'h8000;
LUT4 lut_inst_2720 (
  .F(lut_f_2720),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2720.INIT = 16'h8000;
LUT4 lut_inst_2721 (
  .F(lut_f_2721),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2721.INIT = 16'h8000;
LUT4 lut_inst_2722 (
  .F(lut_f_2722),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2722.INIT = 16'h8000;
LUT4 lut_inst_2723 (
  .F(lut_f_2723),
  .I0(lut_f_2720),
  .I1(lut_f_2721),
  .I2(lut_f_2722),
  .I3(gw_vcc)
);
defparam lut_inst_2723.INIT = 16'h8000;
LUT4 lut_inst_2724 (
  .F(lut_f_2724),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2724.INIT = 16'h8000;
LUT4 lut_inst_2725 (
  .F(lut_f_2725),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2725.INIT = 16'h8000;
LUT4 lut_inst_2726 (
  .F(lut_f_2726),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2726.INIT = 16'h8000;
LUT4 lut_inst_2727 (
  .F(lut_f_2727),
  .I0(lut_f_2724),
  .I1(lut_f_2725),
  .I2(lut_f_2726),
  .I3(gw_vcc)
);
defparam lut_inst_2727.INIT = 16'h8000;
LUT4 lut_inst_2728 (
  .F(lut_f_2728),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2728.INIT = 16'h8000;
LUT4 lut_inst_2729 (
  .F(lut_f_2729),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2729.INIT = 16'h8000;
LUT4 lut_inst_2730 (
  .F(lut_f_2730),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2730.INIT = 16'h8000;
LUT4 lut_inst_2731 (
  .F(lut_f_2731),
  .I0(lut_f_2728),
  .I1(lut_f_2729),
  .I2(lut_f_2730),
  .I3(gw_vcc)
);
defparam lut_inst_2731.INIT = 16'h8000;
LUT4 lut_inst_2732 (
  .F(lut_f_2732),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2732.INIT = 16'h8000;
LUT4 lut_inst_2733 (
  .F(lut_f_2733),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2733.INIT = 16'h8000;
LUT4 lut_inst_2734 (
  .F(lut_f_2734),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2734.INIT = 16'h8000;
LUT4 lut_inst_2735 (
  .F(lut_f_2735),
  .I0(lut_f_2732),
  .I1(lut_f_2733),
  .I2(lut_f_2734),
  .I3(gw_vcc)
);
defparam lut_inst_2735.INIT = 16'h8000;
LUT4 lut_inst_2736 (
  .F(lut_f_2736),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2736.INIT = 16'h8000;
LUT4 lut_inst_2737 (
  .F(lut_f_2737),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2737.INIT = 16'h8000;
LUT4 lut_inst_2738 (
  .F(lut_f_2738),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2738.INIT = 16'h8000;
LUT4 lut_inst_2739 (
  .F(lut_f_2739),
  .I0(lut_f_2736),
  .I1(lut_f_2737),
  .I2(lut_f_2738),
  .I3(gw_vcc)
);
defparam lut_inst_2739.INIT = 16'h8000;
LUT4 lut_inst_2740 (
  .F(lut_f_2740),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2740.INIT = 16'h8000;
LUT4 lut_inst_2741 (
  .F(lut_f_2741),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2741.INIT = 16'h8000;
LUT4 lut_inst_2742 (
  .F(lut_f_2742),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2742.INIT = 16'h8000;
LUT4 lut_inst_2743 (
  .F(lut_f_2743),
  .I0(lut_f_2740),
  .I1(lut_f_2741),
  .I2(lut_f_2742),
  .I3(gw_vcc)
);
defparam lut_inst_2743.INIT = 16'h8000;
LUT4 lut_inst_2744 (
  .F(lut_f_2744),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2744.INIT = 16'h8000;
LUT4 lut_inst_2745 (
  .F(lut_f_2745),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2745.INIT = 16'h8000;
LUT4 lut_inst_2746 (
  .F(lut_f_2746),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2746.INIT = 16'h8000;
LUT4 lut_inst_2747 (
  .F(lut_f_2747),
  .I0(lut_f_2744),
  .I1(lut_f_2745),
  .I2(lut_f_2746),
  .I3(gw_vcc)
);
defparam lut_inst_2747.INIT = 16'h8000;
LUT4 lut_inst_2748 (
  .F(lut_f_2748),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2748.INIT = 16'h8000;
LUT4 lut_inst_2749 (
  .F(lut_f_2749),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2749.INIT = 16'h8000;
LUT4 lut_inst_2750 (
  .F(lut_f_2750),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2750.INIT = 16'h8000;
LUT4 lut_inst_2751 (
  .F(lut_f_2751),
  .I0(lut_f_2748),
  .I1(lut_f_2749),
  .I2(lut_f_2750),
  .I3(gw_vcc)
);
defparam lut_inst_2751.INIT = 16'h8000;
LUT4 lut_inst_2752 (
  .F(lut_f_2752),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2752.INIT = 16'h8000;
LUT4 lut_inst_2753 (
  .F(lut_f_2753),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2753.INIT = 16'h8000;
LUT4 lut_inst_2754 (
  .F(lut_f_2754),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2754.INIT = 16'h8000;
LUT4 lut_inst_2755 (
  .F(lut_f_2755),
  .I0(lut_f_2752),
  .I1(lut_f_2753),
  .I2(lut_f_2754),
  .I3(gw_vcc)
);
defparam lut_inst_2755.INIT = 16'h8000;
LUT4 lut_inst_2756 (
  .F(lut_f_2756),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2756.INIT = 16'h8000;
LUT4 lut_inst_2757 (
  .F(lut_f_2757),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2757.INIT = 16'h8000;
LUT4 lut_inst_2758 (
  .F(lut_f_2758),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2758.INIT = 16'h8000;
LUT4 lut_inst_2759 (
  .F(lut_f_2759),
  .I0(lut_f_2756),
  .I1(lut_f_2757),
  .I2(lut_f_2758),
  .I3(gw_vcc)
);
defparam lut_inst_2759.INIT = 16'h8000;
LUT4 lut_inst_2760 (
  .F(lut_f_2760),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2760.INIT = 16'h8000;
LUT4 lut_inst_2761 (
  .F(lut_f_2761),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2761.INIT = 16'h8000;
LUT4 lut_inst_2762 (
  .F(lut_f_2762),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2762.INIT = 16'h8000;
LUT4 lut_inst_2763 (
  .F(lut_f_2763),
  .I0(lut_f_2760),
  .I1(lut_f_2761),
  .I2(lut_f_2762),
  .I3(gw_vcc)
);
defparam lut_inst_2763.INIT = 16'h8000;
LUT4 lut_inst_2764 (
  .F(lut_f_2764),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2764.INIT = 16'h8000;
LUT4 lut_inst_2765 (
  .F(lut_f_2765),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2765.INIT = 16'h8000;
LUT4 lut_inst_2766 (
  .F(lut_f_2766),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2766.INIT = 16'h8000;
LUT4 lut_inst_2767 (
  .F(lut_f_2767),
  .I0(lut_f_2764),
  .I1(lut_f_2765),
  .I2(lut_f_2766),
  .I3(gw_vcc)
);
defparam lut_inst_2767.INIT = 16'h8000;
LUT4 lut_inst_2768 (
  .F(lut_f_2768),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2768.INIT = 16'h8000;
LUT4 lut_inst_2769 (
  .F(lut_f_2769),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2769.INIT = 16'h8000;
LUT4 lut_inst_2770 (
  .F(lut_f_2770),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2770.INIT = 16'h8000;
LUT4 lut_inst_2771 (
  .F(lut_f_2771),
  .I0(lut_f_2768),
  .I1(lut_f_2769),
  .I2(lut_f_2770),
  .I3(gw_vcc)
);
defparam lut_inst_2771.INIT = 16'h8000;
LUT4 lut_inst_2772 (
  .F(lut_f_2772),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2772.INIT = 16'h8000;
LUT4 lut_inst_2773 (
  .F(lut_f_2773),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2773.INIT = 16'h8000;
LUT4 lut_inst_2774 (
  .F(lut_f_2774),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2774.INIT = 16'h8000;
LUT4 lut_inst_2775 (
  .F(lut_f_2775),
  .I0(lut_f_2772),
  .I1(lut_f_2773),
  .I2(lut_f_2774),
  .I3(gw_vcc)
);
defparam lut_inst_2775.INIT = 16'h8000;
LUT4 lut_inst_2776 (
  .F(lut_f_2776),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2776.INIT = 16'h8000;
LUT4 lut_inst_2777 (
  .F(lut_f_2777),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2777.INIT = 16'h8000;
LUT4 lut_inst_2778 (
  .F(lut_f_2778),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2778.INIT = 16'h8000;
LUT4 lut_inst_2779 (
  .F(lut_f_2779),
  .I0(lut_f_2776),
  .I1(lut_f_2777),
  .I2(lut_f_2778),
  .I3(gw_vcc)
);
defparam lut_inst_2779.INIT = 16'h8000;
LUT4 lut_inst_2780 (
  .F(lut_f_2780),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2780.INIT = 16'h8000;
LUT4 lut_inst_2781 (
  .F(lut_f_2781),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2781.INIT = 16'h8000;
LUT4 lut_inst_2782 (
  .F(lut_f_2782),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2782.INIT = 16'h8000;
LUT4 lut_inst_2783 (
  .F(lut_f_2783),
  .I0(lut_f_2780),
  .I1(lut_f_2781),
  .I2(lut_f_2782),
  .I3(gw_vcc)
);
defparam lut_inst_2783.INIT = 16'h8000;
LUT4 lut_inst_2784 (
  .F(lut_f_2784),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2784.INIT = 16'h8000;
LUT4 lut_inst_2785 (
  .F(lut_f_2785),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2785.INIT = 16'h8000;
LUT4 lut_inst_2786 (
  .F(lut_f_2786),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2786.INIT = 16'h8000;
LUT4 lut_inst_2787 (
  .F(lut_f_2787),
  .I0(lut_f_2784),
  .I1(lut_f_2785),
  .I2(lut_f_2786),
  .I3(gw_vcc)
);
defparam lut_inst_2787.INIT = 16'h8000;
LUT4 lut_inst_2788 (
  .F(lut_f_2788),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2788.INIT = 16'h8000;
LUT4 lut_inst_2789 (
  .F(lut_f_2789),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2789.INIT = 16'h8000;
LUT4 lut_inst_2790 (
  .F(lut_f_2790),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2790.INIT = 16'h8000;
LUT4 lut_inst_2791 (
  .F(lut_f_2791),
  .I0(lut_f_2788),
  .I1(lut_f_2789),
  .I2(lut_f_2790),
  .I3(gw_vcc)
);
defparam lut_inst_2791.INIT = 16'h8000;
LUT4 lut_inst_2792 (
  .F(lut_f_2792),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2792.INIT = 16'h8000;
LUT4 lut_inst_2793 (
  .F(lut_f_2793),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2793.INIT = 16'h8000;
LUT4 lut_inst_2794 (
  .F(lut_f_2794),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2794.INIT = 16'h8000;
LUT4 lut_inst_2795 (
  .F(lut_f_2795),
  .I0(lut_f_2792),
  .I1(lut_f_2793),
  .I2(lut_f_2794),
  .I3(gw_vcc)
);
defparam lut_inst_2795.INIT = 16'h8000;
LUT4 lut_inst_2796 (
  .F(lut_f_2796),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2796.INIT = 16'h8000;
LUT4 lut_inst_2797 (
  .F(lut_f_2797),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2797.INIT = 16'h8000;
LUT4 lut_inst_2798 (
  .F(lut_f_2798),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2798.INIT = 16'h8000;
LUT4 lut_inst_2799 (
  .F(lut_f_2799),
  .I0(lut_f_2796),
  .I1(lut_f_2797),
  .I2(lut_f_2798),
  .I3(gw_vcc)
);
defparam lut_inst_2799.INIT = 16'h8000;
LUT4 lut_inst_2800 (
  .F(lut_f_2800),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2800.INIT = 16'h8000;
LUT4 lut_inst_2801 (
  .F(lut_f_2801),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2801.INIT = 16'h8000;
LUT4 lut_inst_2802 (
  .F(lut_f_2802),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2802.INIT = 16'h8000;
LUT4 lut_inst_2803 (
  .F(lut_f_2803),
  .I0(lut_f_2800),
  .I1(lut_f_2801),
  .I2(lut_f_2802),
  .I3(gw_vcc)
);
defparam lut_inst_2803.INIT = 16'h8000;
LUT4 lut_inst_2804 (
  .F(lut_f_2804),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2804.INIT = 16'h8000;
LUT4 lut_inst_2805 (
  .F(lut_f_2805),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2805.INIT = 16'h8000;
LUT4 lut_inst_2806 (
  .F(lut_f_2806),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2806.INIT = 16'h8000;
LUT4 lut_inst_2807 (
  .F(lut_f_2807),
  .I0(lut_f_2804),
  .I1(lut_f_2805),
  .I2(lut_f_2806),
  .I3(gw_vcc)
);
defparam lut_inst_2807.INIT = 16'h8000;
LUT4 lut_inst_2808 (
  .F(lut_f_2808),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2808.INIT = 16'h8000;
LUT4 lut_inst_2809 (
  .F(lut_f_2809),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2809.INIT = 16'h8000;
LUT4 lut_inst_2810 (
  .F(lut_f_2810),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2810.INIT = 16'h8000;
LUT4 lut_inst_2811 (
  .F(lut_f_2811),
  .I0(lut_f_2808),
  .I1(lut_f_2809),
  .I2(lut_f_2810),
  .I3(gw_vcc)
);
defparam lut_inst_2811.INIT = 16'h8000;
LUT4 lut_inst_2812 (
  .F(lut_f_2812),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2812.INIT = 16'h8000;
LUT4 lut_inst_2813 (
  .F(lut_f_2813),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad10_inv)
);
defparam lut_inst_2813.INIT = 16'h8000;
LUT4 lut_inst_2814 (
  .F(lut_f_2814),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2814.INIT = 16'h8000;
LUT4 lut_inst_2815 (
  .F(lut_f_2815),
  .I0(lut_f_2812),
  .I1(lut_f_2813),
  .I2(lut_f_2814),
  .I3(gw_vcc)
);
defparam lut_inst_2815.INIT = 16'h8000;
LUT4 lut_inst_2816 (
  .F(lut_f_2816),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2816.INIT = 16'h8000;
LUT4 lut_inst_2817 (
  .F(lut_f_2817),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2817.INIT = 16'h8000;
LUT4 lut_inst_2818 (
  .F(lut_f_2818),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2818.INIT = 16'h8000;
LUT4 lut_inst_2819 (
  .F(lut_f_2819),
  .I0(lut_f_2816),
  .I1(lut_f_2817),
  .I2(lut_f_2818),
  .I3(gw_vcc)
);
defparam lut_inst_2819.INIT = 16'h8000;
LUT4 lut_inst_2820 (
  .F(lut_f_2820),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2820.INIT = 16'h8000;
LUT4 lut_inst_2821 (
  .F(lut_f_2821),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2821.INIT = 16'h8000;
LUT4 lut_inst_2822 (
  .F(lut_f_2822),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2822.INIT = 16'h8000;
LUT4 lut_inst_2823 (
  .F(lut_f_2823),
  .I0(lut_f_2820),
  .I1(lut_f_2821),
  .I2(lut_f_2822),
  .I3(gw_vcc)
);
defparam lut_inst_2823.INIT = 16'h8000;
LUT4 lut_inst_2824 (
  .F(lut_f_2824),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2824.INIT = 16'h8000;
LUT4 lut_inst_2825 (
  .F(lut_f_2825),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2825.INIT = 16'h8000;
LUT4 lut_inst_2826 (
  .F(lut_f_2826),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2826.INIT = 16'h8000;
LUT4 lut_inst_2827 (
  .F(lut_f_2827),
  .I0(lut_f_2824),
  .I1(lut_f_2825),
  .I2(lut_f_2826),
  .I3(gw_vcc)
);
defparam lut_inst_2827.INIT = 16'h8000;
LUT4 lut_inst_2828 (
  .F(lut_f_2828),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2828.INIT = 16'h8000;
LUT4 lut_inst_2829 (
  .F(lut_f_2829),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2829.INIT = 16'h8000;
LUT4 lut_inst_2830 (
  .F(lut_f_2830),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2830.INIT = 16'h8000;
LUT4 lut_inst_2831 (
  .F(lut_f_2831),
  .I0(lut_f_2828),
  .I1(lut_f_2829),
  .I2(lut_f_2830),
  .I3(gw_vcc)
);
defparam lut_inst_2831.INIT = 16'h8000;
LUT4 lut_inst_2832 (
  .F(lut_f_2832),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2832.INIT = 16'h8000;
LUT4 lut_inst_2833 (
  .F(lut_f_2833),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2833.INIT = 16'h8000;
LUT4 lut_inst_2834 (
  .F(lut_f_2834),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2834.INIT = 16'h8000;
LUT4 lut_inst_2835 (
  .F(lut_f_2835),
  .I0(lut_f_2832),
  .I1(lut_f_2833),
  .I2(lut_f_2834),
  .I3(gw_vcc)
);
defparam lut_inst_2835.INIT = 16'h8000;
LUT4 lut_inst_2836 (
  .F(lut_f_2836),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2836.INIT = 16'h8000;
LUT4 lut_inst_2837 (
  .F(lut_f_2837),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2837.INIT = 16'h8000;
LUT4 lut_inst_2838 (
  .F(lut_f_2838),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2838.INIT = 16'h8000;
LUT4 lut_inst_2839 (
  .F(lut_f_2839),
  .I0(lut_f_2836),
  .I1(lut_f_2837),
  .I2(lut_f_2838),
  .I3(gw_vcc)
);
defparam lut_inst_2839.INIT = 16'h8000;
LUT4 lut_inst_2840 (
  .F(lut_f_2840),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2840.INIT = 16'h8000;
LUT4 lut_inst_2841 (
  .F(lut_f_2841),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2841.INIT = 16'h8000;
LUT4 lut_inst_2842 (
  .F(lut_f_2842),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2842.INIT = 16'h8000;
LUT4 lut_inst_2843 (
  .F(lut_f_2843),
  .I0(lut_f_2840),
  .I1(lut_f_2841),
  .I2(lut_f_2842),
  .I3(gw_vcc)
);
defparam lut_inst_2843.INIT = 16'h8000;
LUT4 lut_inst_2844 (
  .F(lut_f_2844),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2844.INIT = 16'h8000;
LUT4 lut_inst_2845 (
  .F(lut_f_2845),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2845.INIT = 16'h8000;
LUT4 lut_inst_2846 (
  .F(lut_f_2846),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2846.INIT = 16'h8000;
LUT4 lut_inst_2847 (
  .F(lut_f_2847),
  .I0(lut_f_2844),
  .I1(lut_f_2845),
  .I2(lut_f_2846),
  .I3(gw_vcc)
);
defparam lut_inst_2847.INIT = 16'h8000;
LUT4 lut_inst_2848 (
  .F(lut_f_2848),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2848.INIT = 16'h8000;
LUT4 lut_inst_2849 (
  .F(lut_f_2849),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2849.INIT = 16'h8000;
LUT4 lut_inst_2850 (
  .F(lut_f_2850),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2850.INIT = 16'h8000;
LUT4 lut_inst_2851 (
  .F(lut_f_2851),
  .I0(lut_f_2848),
  .I1(lut_f_2849),
  .I2(lut_f_2850),
  .I3(gw_vcc)
);
defparam lut_inst_2851.INIT = 16'h8000;
LUT4 lut_inst_2852 (
  .F(lut_f_2852),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2852.INIT = 16'h8000;
LUT4 lut_inst_2853 (
  .F(lut_f_2853),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2853.INIT = 16'h8000;
LUT4 lut_inst_2854 (
  .F(lut_f_2854),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2854.INIT = 16'h8000;
LUT4 lut_inst_2855 (
  .F(lut_f_2855),
  .I0(lut_f_2852),
  .I1(lut_f_2853),
  .I2(lut_f_2854),
  .I3(gw_vcc)
);
defparam lut_inst_2855.INIT = 16'h8000;
LUT4 lut_inst_2856 (
  .F(lut_f_2856),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2856.INIT = 16'h8000;
LUT4 lut_inst_2857 (
  .F(lut_f_2857),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2857.INIT = 16'h8000;
LUT4 lut_inst_2858 (
  .F(lut_f_2858),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2858.INIT = 16'h8000;
LUT4 lut_inst_2859 (
  .F(lut_f_2859),
  .I0(lut_f_2856),
  .I1(lut_f_2857),
  .I2(lut_f_2858),
  .I3(gw_vcc)
);
defparam lut_inst_2859.INIT = 16'h8000;
LUT4 lut_inst_2860 (
  .F(lut_f_2860),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2860.INIT = 16'h8000;
LUT4 lut_inst_2861 (
  .F(lut_f_2861),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2861.INIT = 16'h8000;
LUT4 lut_inst_2862 (
  .F(lut_f_2862),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2862.INIT = 16'h8000;
LUT4 lut_inst_2863 (
  .F(lut_f_2863),
  .I0(lut_f_2860),
  .I1(lut_f_2861),
  .I2(lut_f_2862),
  .I3(gw_vcc)
);
defparam lut_inst_2863.INIT = 16'h8000;
LUT4 lut_inst_2864 (
  .F(lut_f_2864),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2864.INIT = 16'h8000;
LUT4 lut_inst_2865 (
  .F(lut_f_2865),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2865.INIT = 16'h8000;
LUT4 lut_inst_2866 (
  .F(lut_f_2866),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2866.INIT = 16'h8000;
LUT4 lut_inst_2867 (
  .F(lut_f_2867),
  .I0(lut_f_2864),
  .I1(lut_f_2865),
  .I2(lut_f_2866),
  .I3(gw_vcc)
);
defparam lut_inst_2867.INIT = 16'h8000;
LUT4 lut_inst_2868 (
  .F(lut_f_2868),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2868.INIT = 16'h8000;
LUT4 lut_inst_2869 (
  .F(lut_f_2869),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2869.INIT = 16'h8000;
LUT4 lut_inst_2870 (
  .F(lut_f_2870),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2870.INIT = 16'h8000;
LUT4 lut_inst_2871 (
  .F(lut_f_2871),
  .I0(lut_f_2868),
  .I1(lut_f_2869),
  .I2(lut_f_2870),
  .I3(gw_vcc)
);
defparam lut_inst_2871.INIT = 16'h8000;
LUT4 lut_inst_2872 (
  .F(lut_f_2872),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2872.INIT = 16'h8000;
LUT4 lut_inst_2873 (
  .F(lut_f_2873),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2873.INIT = 16'h8000;
LUT4 lut_inst_2874 (
  .F(lut_f_2874),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2874.INIT = 16'h8000;
LUT4 lut_inst_2875 (
  .F(lut_f_2875),
  .I0(lut_f_2872),
  .I1(lut_f_2873),
  .I2(lut_f_2874),
  .I3(gw_vcc)
);
defparam lut_inst_2875.INIT = 16'h8000;
LUT4 lut_inst_2876 (
  .F(lut_f_2876),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2876.INIT = 16'h8000;
LUT4 lut_inst_2877 (
  .F(lut_f_2877),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2877.INIT = 16'h8000;
LUT4 lut_inst_2878 (
  .F(lut_f_2878),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2878.INIT = 16'h8000;
LUT4 lut_inst_2879 (
  .F(lut_f_2879),
  .I0(lut_f_2876),
  .I1(lut_f_2877),
  .I2(lut_f_2878),
  .I3(gw_vcc)
);
defparam lut_inst_2879.INIT = 16'h8000;
LUT4 lut_inst_2880 (
  .F(lut_f_2880),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2880.INIT = 16'h8000;
LUT4 lut_inst_2881 (
  .F(lut_f_2881),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2881.INIT = 16'h8000;
LUT4 lut_inst_2882 (
  .F(lut_f_2882),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2882.INIT = 16'h8000;
LUT4 lut_inst_2883 (
  .F(lut_f_2883),
  .I0(lut_f_2880),
  .I1(lut_f_2881),
  .I2(lut_f_2882),
  .I3(gw_vcc)
);
defparam lut_inst_2883.INIT = 16'h8000;
LUT4 lut_inst_2884 (
  .F(lut_f_2884),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2884.INIT = 16'h8000;
LUT4 lut_inst_2885 (
  .F(lut_f_2885),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2885.INIT = 16'h8000;
LUT4 lut_inst_2886 (
  .F(lut_f_2886),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2886.INIT = 16'h8000;
LUT4 lut_inst_2887 (
  .F(lut_f_2887),
  .I0(lut_f_2884),
  .I1(lut_f_2885),
  .I2(lut_f_2886),
  .I3(gw_vcc)
);
defparam lut_inst_2887.INIT = 16'h8000;
LUT4 lut_inst_2888 (
  .F(lut_f_2888),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2888.INIT = 16'h8000;
LUT4 lut_inst_2889 (
  .F(lut_f_2889),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2889.INIT = 16'h8000;
LUT4 lut_inst_2890 (
  .F(lut_f_2890),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2890.INIT = 16'h8000;
LUT4 lut_inst_2891 (
  .F(lut_f_2891),
  .I0(lut_f_2888),
  .I1(lut_f_2889),
  .I2(lut_f_2890),
  .I3(gw_vcc)
);
defparam lut_inst_2891.INIT = 16'h8000;
LUT4 lut_inst_2892 (
  .F(lut_f_2892),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2892.INIT = 16'h8000;
LUT4 lut_inst_2893 (
  .F(lut_f_2893),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2893.INIT = 16'h8000;
LUT4 lut_inst_2894 (
  .F(lut_f_2894),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2894.INIT = 16'h8000;
LUT4 lut_inst_2895 (
  .F(lut_f_2895),
  .I0(lut_f_2892),
  .I1(lut_f_2893),
  .I2(lut_f_2894),
  .I3(gw_vcc)
);
defparam lut_inst_2895.INIT = 16'h8000;
LUT4 lut_inst_2896 (
  .F(lut_f_2896),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2896.INIT = 16'h8000;
LUT4 lut_inst_2897 (
  .F(lut_f_2897),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2897.INIT = 16'h8000;
LUT4 lut_inst_2898 (
  .F(lut_f_2898),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2898.INIT = 16'h8000;
LUT4 lut_inst_2899 (
  .F(lut_f_2899),
  .I0(lut_f_2896),
  .I1(lut_f_2897),
  .I2(lut_f_2898),
  .I3(gw_vcc)
);
defparam lut_inst_2899.INIT = 16'h8000;
LUT4 lut_inst_2900 (
  .F(lut_f_2900),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2900.INIT = 16'h8000;
LUT4 lut_inst_2901 (
  .F(lut_f_2901),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2901.INIT = 16'h8000;
LUT4 lut_inst_2902 (
  .F(lut_f_2902),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2902.INIT = 16'h8000;
LUT4 lut_inst_2903 (
  .F(lut_f_2903),
  .I0(lut_f_2900),
  .I1(lut_f_2901),
  .I2(lut_f_2902),
  .I3(gw_vcc)
);
defparam lut_inst_2903.INIT = 16'h8000;
LUT4 lut_inst_2904 (
  .F(lut_f_2904),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2904.INIT = 16'h8000;
LUT4 lut_inst_2905 (
  .F(lut_f_2905),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2905.INIT = 16'h8000;
LUT4 lut_inst_2906 (
  .F(lut_f_2906),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2906.INIT = 16'h8000;
LUT4 lut_inst_2907 (
  .F(lut_f_2907),
  .I0(lut_f_2904),
  .I1(lut_f_2905),
  .I2(lut_f_2906),
  .I3(gw_vcc)
);
defparam lut_inst_2907.INIT = 16'h8000;
LUT4 lut_inst_2908 (
  .F(lut_f_2908),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2908.INIT = 16'h8000;
LUT4 lut_inst_2909 (
  .F(lut_f_2909),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2909.INIT = 16'h8000;
LUT4 lut_inst_2910 (
  .F(lut_f_2910),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2910.INIT = 16'h8000;
LUT4 lut_inst_2911 (
  .F(lut_f_2911),
  .I0(lut_f_2908),
  .I1(lut_f_2909),
  .I2(lut_f_2910),
  .I3(gw_vcc)
);
defparam lut_inst_2911.INIT = 16'h8000;
LUT4 lut_inst_2912 (
  .F(lut_f_2912),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2912.INIT = 16'h8000;
LUT4 lut_inst_2913 (
  .F(lut_f_2913),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2913.INIT = 16'h8000;
LUT4 lut_inst_2914 (
  .F(lut_f_2914),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2914.INIT = 16'h8000;
LUT4 lut_inst_2915 (
  .F(lut_f_2915),
  .I0(lut_f_2912),
  .I1(lut_f_2913),
  .I2(lut_f_2914),
  .I3(gw_vcc)
);
defparam lut_inst_2915.INIT = 16'h8000;
LUT4 lut_inst_2916 (
  .F(lut_f_2916),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2916.INIT = 16'h8000;
LUT4 lut_inst_2917 (
  .F(lut_f_2917),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2917.INIT = 16'h8000;
LUT4 lut_inst_2918 (
  .F(lut_f_2918),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2918.INIT = 16'h8000;
LUT4 lut_inst_2919 (
  .F(lut_f_2919),
  .I0(lut_f_2916),
  .I1(lut_f_2917),
  .I2(lut_f_2918),
  .I3(gw_vcc)
);
defparam lut_inst_2919.INIT = 16'h8000;
LUT4 lut_inst_2920 (
  .F(lut_f_2920),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2920.INIT = 16'h8000;
LUT4 lut_inst_2921 (
  .F(lut_f_2921),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2921.INIT = 16'h8000;
LUT4 lut_inst_2922 (
  .F(lut_f_2922),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2922.INIT = 16'h8000;
LUT4 lut_inst_2923 (
  .F(lut_f_2923),
  .I0(lut_f_2920),
  .I1(lut_f_2921),
  .I2(lut_f_2922),
  .I3(gw_vcc)
);
defparam lut_inst_2923.INIT = 16'h8000;
LUT4 lut_inst_2924 (
  .F(lut_f_2924),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2924.INIT = 16'h8000;
LUT4 lut_inst_2925 (
  .F(lut_f_2925),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2925.INIT = 16'h8000;
LUT4 lut_inst_2926 (
  .F(lut_f_2926),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2926.INIT = 16'h8000;
LUT4 lut_inst_2927 (
  .F(lut_f_2927),
  .I0(lut_f_2924),
  .I1(lut_f_2925),
  .I2(lut_f_2926),
  .I3(gw_vcc)
);
defparam lut_inst_2927.INIT = 16'h8000;
LUT4 lut_inst_2928 (
  .F(lut_f_2928),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2928.INIT = 16'h8000;
LUT4 lut_inst_2929 (
  .F(lut_f_2929),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2929.INIT = 16'h8000;
LUT4 lut_inst_2930 (
  .F(lut_f_2930),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2930.INIT = 16'h8000;
LUT4 lut_inst_2931 (
  .F(lut_f_2931),
  .I0(lut_f_2928),
  .I1(lut_f_2929),
  .I2(lut_f_2930),
  .I3(gw_vcc)
);
defparam lut_inst_2931.INIT = 16'h8000;
LUT4 lut_inst_2932 (
  .F(lut_f_2932),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2932.INIT = 16'h8000;
LUT4 lut_inst_2933 (
  .F(lut_f_2933),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2933.INIT = 16'h8000;
LUT4 lut_inst_2934 (
  .F(lut_f_2934),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2934.INIT = 16'h8000;
LUT4 lut_inst_2935 (
  .F(lut_f_2935),
  .I0(lut_f_2932),
  .I1(lut_f_2933),
  .I2(lut_f_2934),
  .I3(gw_vcc)
);
defparam lut_inst_2935.INIT = 16'h8000;
LUT4 lut_inst_2936 (
  .F(lut_f_2936),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2936.INIT = 16'h8000;
LUT4 lut_inst_2937 (
  .F(lut_f_2937),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2937.INIT = 16'h8000;
LUT4 lut_inst_2938 (
  .F(lut_f_2938),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2938.INIT = 16'h8000;
LUT4 lut_inst_2939 (
  .F(lut_f_2939),
  .I0(lut_f_2936),
  .I1(lut_f_2937),
  .I2(lut_f_2938),
  .I3(gw_vcc)
);
defparam lut_inst_2939.INIT = 16'h8000;
LUT4 lut_inst_2940 (
  .F(lut_f_2940),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2940.INIT = 16'h8000;
LUT4 lut_inst_2941 (
  .F(lut_f_2941),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad[10])
);
defparam lut_inst_2941.INIT = 16'h8000;
LUT4 lut_inst_2942 (
  .F(lut_f_2942),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2942.INIT = 16'h8000;
LUT4 lut_inst_2943 (
  .F(lut_f_2943),
  .I0(lut_f_2940),
  .I1(lut_f_2941),
  .I2(lut_f_2942),
  .I3(gw_vcc)
);
defparam lut_inst_2943.INIT = 16'h8000;
LUT4 lut_inst_2944 (
  .F(lut_f_2944),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2944.INIT = 16'h8000;
LUT4 lut_inst_2945 (
  .F(lut_f_2945),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2945.INIT = 16'h8000;
LUT4 lut_inst_2946 (
  .F(lut_f_2946),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2946.INIT = 16'h8000;
LUT4 lut_inst_2947 (
  .F(lut_f_2947),
  .I0(lut_f_2944),
  .I1(lut_f_2945),
  .I2(lut_f_2946),
  .I3(gw_vcc)
);
defparam lut_inst_2947.INIT = 16'h8000;
LUT4 lut_inst_2948 (
  .F(lut_f_2948),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2948.INIT = 16'h8000;
LUT4 lut_inst_2949 (
  .F(lut_f_2949),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2949.INIT = 16'h8000;
LUT4 lut_inst_2950 (
  .F(lut_f_2950),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2950.INIT = 16'h8000;
LUT4 lut_inst_2951 (
  .F(lut_f_2951),
  .I0(lut_f_2948),
  .I1(lut_f_2949),
  .I2(lut_f_2950),
  .I3(gw_vcc)
);
defparam lut_inst_2951.INIT = 16'h8000;
LUT4 lut_inst_2952 (
  .F(lut_f_2952),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2952.INIT = 16'h8000;
LUT4 lut_inst_2953 (
  .F(lut_f_2953),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2953.INIT = 16'h8000;
LUT4 lut_inst_2954 (
  .F(lut_f_2954),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2954.INIT = 16'h8000;
LUT4 lut_inst_2955 (
  .F(lut_f_2955),
  .I0(lut_f_2952),
  .I1(lut_f_2953),
  .I2(lut_f_2954),
  .I3(gw_vcc)
);
defparam lut_inst_2955.INIT = 16'h8000;
LUT4 lut_inst_2956 (
  .F(lut_f_2956),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2956.INIT = 16'h8000;
LUT4 lut_inst_2957 (
  .F(lut_f_2957),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2957.INIT = 16'h8000;
LUT4 lut_inst_2958 (
  .F(lut_f_2958),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2958.INIT = 16'h8000;
LUT4 lut_inst_2959 (
  .F(lut_f_2959),
  .I0(lut_f_2956),
  .I1(lut_f_2957),
  .I2(lut_f_2958),
  .I3(gw_vcc)
);
defparam lut_inst_2959.INIT = 16'h8000;
LUT4 lut_inst_2960 (
  .F(lut_f_2960),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2960.INIT = 16'h8000;
LUT4 lut_inst_2961 (
  .F(lut_f_2961),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2961.INIT = 16'h8000;
LUT4 lut_inst_2962 (
  .F(lut_f_2962),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2962.INIT = 16'h8000;
LUT4 lut_inst_2963 (
  .F(lut_f_2963),
  .I0(lut_f_2960),
  .I1(lut_f_2961),
  .I2(lut_f_2962),
  .I3(gw_vcc)
);
defparam lut_inst_2963.INIT = 16'h8000;
LUT4 lut_inst_2964 (
  .F(lut_f_2964),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2964.INIT = 16'h8000;
LUT4 lut_inst_2965 (
  .F(lut_f_2965),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2965.INIT = 16'h8000;
LUT4 lut_inst_2966 (
  .F(lut_f_2966),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2966.INIT = 16'h8000;
LUT4 lut_inst_2967 (
  .F(lut_f_2967),
  .I0(lut_f_2964),
  .I1(lut_f_2965),
  .I2(lut_f_2966),
  .I3(gw_vcc)
);
defparam lut_inst_2967.INIT = 16'h8000;
LUT4 lut_inst_2968 (
  .F(lut_f_2968),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2968.INIT = 16'h8000;
LUT4 lut_inst_2969 (
  .F(lut_f_2969),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2969.INIT = 16'h8000;
LUT4 lut_inst_2970 (
  .F(lut_f_2970),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2970.INIT = 16'h8000;
LUT4 lut_inst_2971 (
  .F(lut_f_2971),
  .I0(lut_f_2968),
  .I1(lut_f_2969),
  .I2(lut_f_2970),
  .I3(gw_vcc)
);
defparam lut_inst_2971.INIT = 16'h8000;
LUT4 lut_inst_2972 (
  .F(lut_f_2972),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_2972.INIT = 16'h8000;
LUT4 lut_inst_2973 (
  .F(lut_f_2973),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2973.INIT = 16'h8000;
LUT4 lut_inst_2974 (
  .F(lut_f_2974),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2974.INIT = 16'h8000;
LUT4 lut_inst_2975 (
  .F(lut_f_2975),
  .I0(lut_f_2972),
  .I1(lut_f_2973),
  .I2(lut_f_2974),
  .I3(gw_vcc)
);
defparam lut_inst_2975.INIT = 16'h8000;
LUT4 lut_inst_2976 (
  .F(lut_f_2976),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2976.INIT = 16'h8000;
LUT4 lut_inst_2977 (
  .F(lut_f_2977),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2977.INIT = 16'h8000;
LUT4 lut_inst_2978 (
  .F(lut_f_2978),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2978.INIT = 16'h8000;
LUT4 lut_inst_2979 (
  .F(lut_f_2979),
  .I0(lut_f_2976),
  .I1(lut_f_2977),
  .I2(lut_f_2978),
  .I3(gw_vcc)
);
defparam lut_inst_2979.INIT = 16'h8000;
LUT4 lut_inst_2980 (
  .F(lut_f_2980),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_2980.INIT = 16'h8000;
LUT4 lut_inst_2981 (
  .F(lut_f_2981),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2981.INIT = 16'h8000;
LUT4 lut_inst_2982 (
  .F(lut_f_2982),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2982.INIT = 16'h8000;
LUT4 lut_inst_2983 (
  .F(lut_f_2983),
  .I0(lut_f_2980),
  .I1(lut_f_2981),
  .I2(lut_f_2982),
  .I3(gw_vcc)
);
defparam lut_inst_2983.INIT = 16'h8000;
LUT4 lut_inst_2984 (
  .F(lut_f_2984),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2984.INIT = 16'h8000;
LUT4 lut_inst_2985 (
  .F(lut_f_2985),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2985.INIT = 16'h8000;
LUT4 lut_inst_2986 (
  .F(lut_f_2986),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2986.INIT = 16'h8000;
LUT4 lut_inst_2987 (
  .F(lut_f_2987),
  .I0(lut_f_2984),
  .I1(lut_f_2985),
  .I2(lut_f_2986),
  .I3(gw_vcc)
);
defparam lut_inst_2987.INIT = 16'h8000;
LUT4 lut_inst_2988 (
  .F(lut_f_2988),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_2988.INIT = 16'h8000;
LUT4 lut_inst_2989 (
  .F(lut_f_2989),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2989.INIT = 16'h8000;
LUT4 lut_inst_2990 (
  .F(lut_f_2990),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2990.INIT = 16'h8000;
LUT4 lut_inst_2991 (
  .F(lut_f_2991),
  .I0(lut_f_2988),
  .I1(lut_f_2989),
  .I2(lut_f_2990),
  .I3(gw_vcc)
);
defparam lut_inst_2991.INIT = 16'h8000;
LUT4 lut_inst_2992 (
  .F(lut_f_2992),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2992.INIT = 16'h8000;
LUT4 lut_inst_2993 (
  .F(lut_f_2993),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2993.INIT = 16'h8000;
LUT4 lut_inst_2994 (
  .F(lut_f_2994),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2994.INIT = 16'h8000;
LUT4 lut_inst_2995 (
  .F(lut_f_2995),
  .I0(lut_f_2992),
  .I1(lut_f_2993),
  .I2(lut_f_2994),
  .I3(gw_vcc)
);
defparam lut_inst_2995.INIT = 16'h8000;
LUT4 lut_inst_2996 (
  .F(lut_f_2996),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_2996.INIT = 16'h8000;
LUT4 lut_inst_2997 (
  .F(lut_f_2997),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_2997.INIT = 16'h8000;
LUT4 lut_inst_2998 (
  .F(lut_f_2998),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_2998.INIT = 16'h8000;
LUT4 lut_inst_2999 (
  .F(lut_f_2999),
  .I0(lut_f_2996),
  .I1(lut_f_2997),
  .I2(lut_f_2998),
  .I3(gw_vcc)
);
defparam lut_inst_2999.INIT = 16'h8000;
LUT4 lut_inst_3000 (
  .F(lut_f_3000),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3000.INIT = 16'h8000;
LUT4 lut_inst_3001 (
  .F(lut_f_3001),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3001.INIT = 16'h8000;
LUT4 lut_inst_3002 (
  .F(lut_f_3002),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3002.INIT = 16'h8000;
LUT4 lut_inst_3003 (
  .F(lut_f_3003),
  .I0(lut_f_3000),
  .I1(lut_f_3001),
  .I2(lut_f_3002),
  .I3(gw_vcc)
);
defparam lut_inst_3003.INIT = 16'h8000;
LUT4 lut_inst_3004 (
  .F(lut_f_3004),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3004.INIT = 16'h8000;
LUT4 lut_inst_3005 (
  .F(lut_f_3005),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3005.INIT = 16'h8000;
LUT4 lut_inst_3006 (
  .F(lut_f_3006),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3006.INIT = 16'h8000;
LUT4 lut_inst_3007 (
  .F(lut_f_3007),
  .I0(lut_f_3004),
  .I1(lut_f_3005),
  .I2(lut_f_3006),
  .I3(gw_vcc)
);
defparam lut_inst_3007.INIT = 16'h8000;
LUT4 lut_inst_3008 (
  .F(lut_f_3008),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_3008.INIT = 16'h8000;
LUT4 lut_inst_3009 (
  .F(lut_f_3009),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3009.INIT = 16'h8000;
LUT4 lut_inst_3010 (
  .F(lut_f_3010),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3010.INIT = 16'h8000;
LUT4 lut_inst_3011 (
  .F(lut_f_3011),
  .I0(lut_f_3008),
  .I1(lut_f_3009),
  .I2(lut_f_3010),
  .I3(gw_vcc)
);
defparam lut_inst_3011.INIT = 16'h8000;
LUT4 lut_inst_3012 (
  .F(lut_f_3012),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_3012.INIT = 16'h8000;
LUT4 lut_inst_3013 (
  .F(lut_f_3013),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3013.INIT = 16'h8000;
LUT4 lut_inst_3014 (
  .F(lut_f_3014),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3014.INIT = 16'h8000;
LUT4 lut_inst_3015 (
  .F(lut_f_3015),
  .I0(lut_f_3012),
  .I1(lut_f_3013),
  .I2(lut_f_3014),
  .I3(gw_vcc)
);
defparam lut_inst_3015.INIT = 16'h8000;
LUT4 lut_inst_3016 (
  .F(lut_f_3016),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_3016.INIT = 16'h8000;
LUT4 lut_inst_3017 (
  .F(lut_f_3017),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3017.INIT = 16'h8000;
LUT4 lut_inst_3018 (
  .F(lut_f_3018),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3018.INIT = 16'h8000;
LUT4 lut_inst_3019 (
  .F(lut_f_3019),
  .I0(lut_f_3016),
  .I1(lut_f_3017),
  .I2(lut_f_3018),
  .I3(gw_vcc)
);
defparam lut_inst_3019.INIT = 16'h8000;
LUT4 lut_inst_3020 (
  .F(lut_f_3020),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_3020.INIT = 16'h8000;
LUT4 lut_inst_3021 (
  .F(lut_f_3021),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3021.INIT = 16'h8000;
LUT4 lut_inst_3022 (
  .F(lut_f_3022),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3022.INIT = 16'h8000;
LUT4 lut_inst_3023 (
  .F(lut_f_3023),
  .I0(lut_f_3020),
  .I1(lut_f_3021),
  .I2(lut_f_3022),
  .I3(gw_vcc)
);
defparam lut_inst_3023.INIT = 16'h8000;
LUT4 lut_inst_3024 (
  .F(lut_f_3024),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_3024.INIT = 16'h8000;
LUT4 lut_inst_3025 (
  .F(lut_f_3025),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3025.INIT = 16'h8000;
LUT4 lut_inst_3026 (
  .F(lut_f_3026),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3026.INIT = 16'h8000;
LUT4 lut_inst_3027 (
  .F(lut_f_3027),
  .I0(lut_f_3024),
  .I1(lut_f_3025),
  .I2(lut_f_3026),
  .I3(gw_vcc)
);
defparam lut_inst_3027.INIT = 16'h8000;
LUT4 lut_inst_3028 (
  .F(lut_f_3028),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_3028.INIT = 16'h8000;
LUT4 lut_inst_3029 (
  .F(lut_f_3029),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3029.INIT = 16'h8000;
LUT4 lut_inst_3030 (
  .F(lut_f_3030),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3030.INIT = 16'h8000;
LUT4 lut_inst_3031 (
  .F(lut_f_3031),
  .I0(lut_f_3028),
  .I1(lut_f_3029),
  .I2(lut_f_3030),
  .I3(gw_vcc)
);
defparam lut_inst_3031.INIT = 16'h8000;
LUT4 lut_inst_3032 (
  .F(lut_f_3032),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3032.INIT = 16'h8000;
LUT4 lut_inst_3033 (
  .F(lut_f_3033),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3033.INIT = 16'h8000;
LUT4 lut_inst_3034 (
  .F(lut_f_3034),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3034.INIT = 16'h8000;
LUT4 lut_inst_3035 (
  .F(lut_f_3035),
  .I0(lut_f_3032),
  .I1(lut_f_3033),
  .I2(lut_f_3034),
  .I3(gw_vcc)
);
defparam lut_inst_3035.INIT = 16'h8000;
LUT4 lut_inst_3036 (
  .F(lut_f_3036),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3036.INIT = 16'h8000;
LUT4 lut_inst_3037 (
  .F(lut_f_3037),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3037.INIT = 16'h8000;
LUT4 lut_inst_3038 (
  .F(lut_f_3038),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3038.INIT = 16'h8000;
LUT4 lut_inst_3039 (
  .F(lut_f_3039),
  .I0(lut_f_3036),
  .I1(lut_f_3037),
  .I2(lut_f_3038),
  .I3(gw_vcc)
);
defparam lut_inst_3039.INIT = 16'h8000;
LUT4 lut_inst_3040 (
  .F(lut_f_3040),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_3040.INIT = 16'h8000;
LUT4 lut_inst_3041 (
  .F(lut_f_3041),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3041.INIT = 16'h8000;
LUT4 lut_inst_3042 (
  .F(lut_f_3042),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3042.INIT = 16'h8000;
LUT4 lut_inst_3043 (
  .F(lut_f_3043),
  .I0(lut_f_3040),
  .I1(lut_f_3041),
  .I2(lut_f_3042),
  .I3(gw_vcc)
);
defparam lut_inst_3043.INIT = 16'h8000;
LUT4 lut_inst_3044 (
  .F(lut_f_3044),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_3044.INIT = 16'h8000;
LUT4 lut_inst_3045 (
  .F(lut_f_3045),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3045.INIT = 16'h8000;
LUT4 lut_inst_3046 (
  .F(lut_f_3046),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3046.INIT = 16'h8000;
LUT4 lut_inst_3047 (
  .F(lut_f_3047),
  .I0(lut_f_3044),
  .I1(lut_f_3045),
  .I2(lut_f_3046),
  .I3(gw_vcc)
);
defparam lut_inst_3047.INIT = 16'h8000;
LUT4 lut_inst_3048 (
  .F(lut_f_3048),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_3048.INIT = 16'h8000;
LUT4 lut_inst_3049 (
  .F(lut_f_3049),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3049.INIT = 16'h8000;
LUT4 lut_inst_3050 (
  .F(lut_f_3050),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3050.INIT = 16'h8000;
LUT4 lut_inst_3051 (
  .F(lut_f_3051),
  .I0(lut_f_3048),
  .I1(lut_f_3049),
  .I2(lut_f_3050),
  .I3(gw_vcc)
);
defparam lut_inst_3051.INIT = 16'h8000;
LUT4 lut_inst_3052 (
  .F(lut_f_3052),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_3052.INIT = 16'h8000;
LUT4 lut_inst_3053 (
  .F(lut_f_3053),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3053.INIT = 16'h8000;
LUT4 lut_inst_3054 (
  .F(lut_f_3054),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3054.INIT = 16'h8000;
LUT4 lut_inst_3055 (
  .F(lut_f_3055),
  .I0(lut_f_3052),
  .I1(lut_f_3053),
  .I2(lut_f_3054),
  .I3(gw_vcc)
);
defparam lut_inst_3055.INIT = 16'h8000;
LUT4 lut_inst_3056 (
  .F(lut_f_3056),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_3056.INIT = 16'h8000;
LUT4 lut_inst_3057 (
  .F(lut_f_3057),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3057.INIT = 16'h8000;
LUT4 lut_inst_3058 (
  .F(lut_f_3058),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3058.INIT = 16'h8000;
LUT4 lut_inst_3059 (
  .F(lut_f_3059),
  .I0(lut_f_3056),
  .I1(lut_f_3057),
  .I2(lut_f_3058),
  .I3(gw_vcc)
);
defparam lut_inst_3059.INIT = 16'h8000;
LUT4 lut_inst_3060 (
  .F(lut_f_3060),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_3060.INIT = 16'h8000;
LUT4 lut_inst_3061 (
  .F(lut_f_3061),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3061.INIT = 16'h8000;
LUT4 lut_inst_3062 (
  .F(lut_f_3062),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3062.INIT = 16'h8000;
LUT4 lut_inst_3063 (
  .F(lut_f_3063),
  .I0(lut_f_3060),
  .I1(lut_f_3061),
  .I2(lut_f_3062),
  .I3(gw_vcc)
);
defparam lut_inst_3063.INIT = 16'h8000;
LUT4 lut_inst_3064 (
  .F(lut_f_3064),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3064.INIT = 16'h8000;
LUT4 lut_inst_3065 (
  .F(lut_f_3065),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3065.INIT = 16'h8000;
LUT4 lut_inst_3066 (
  .F(lut_f_3066),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3066.INIT = 16'h8000;
LUT4 lut_inst_3067 (
  .F(lut_f_3067),
  .I0(lut_f_3064),
  .I1(lut_f_3065),
  .I2(lut_f_3066),
  .I3(gw_vcc)
);
defparam lut_inst_3067.INIT = 16'h8000;
LUT4 lut_inst_3068 (
  .F(lut_f_3068),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3068.INIT = 16'h8000;
LUT4 lut_inst_3069 (
  .F(lut_f_3069),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad[9]),
  .I3(ad[10])
);
defparam lut_inst_3069.INIT = 16'h8000;
LUT4 lut_inst_3070 (
  .F(lut_f_3070),
  .I0(ad[11]),
  .I1(ad12_inv),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3070.INIT = 16'h8000;
LUT4 lut_inst_3071 (
  .F(lut_f_3071),
  .I0(lut_f_3068),
  .I1(lut_f_3069),
  .I2(lut_f_3070),
  .I3(gw_vcc)
);
defparam lut_inst_3071.INIT = 16'h8000;
LUT4 lut_inst_3072 (
  .F(lut_f_3072),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_3072.INIT = 16'h8000;
LUT4 lut_inst_3073 (
  .F(lut_f_3073),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3073.INIT = 16'h8000;
LUT4 lut_inst_3074 (
  .F(lut_f_3074),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3074.INIT = 16'h8000;
LUT4 lut_inst_3075 (
  .F(lut_f_3075),
  .I0(lut_f_3072),
  .I1(lut_f_3073),
  .I2(lut_f_3074),
  .I3(gw_vcc)
);
defparam lut_inst_3075.INIT = 16'h8000;
LUT4 lut_inst_3076 (
  .F(lut_f_3076),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_3076.INIT = 16'h8000;
LUT4 lut_inst_3077 (
  .F(lut_f_3077),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3077.INIT = 16'h8000;
LUT4 lut_inst_3078 (
  .F(lut_f_3078),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3078.INIT = 16'h8000;
LUT4 lut_inst_3079 (
  .F(lut_f_3079),
  .I0(lut_f_3076),
  .I1(lut_f_3077),
  .I2(lut_f_3078),
  .I3(gw_vcc)
);
defparam lut_inst_3079.INIT = 16'h8000;
LUT4 lut_inst_3080 (
  .F(lut_f_3080),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_3080.INIT = 16'h8000;
LUT4 lut_inst_3081 (
  .F(lut_f_3081),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3081.INIT = 16'h8000;
LUT4 lut_inst_3082 (
  .F(lut_f_3082),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3082.INIT = 16'h8000;
LUT4 lut_inst_3083 (
  .F(lut_f_3083),
  .I0(lut_f_3080),
  .I1(lut_f_3081),
  .I2(lut_f_3082),
  .I3(gw_vcc)
);
defparam lut_inst_3083.INIT = 16'h8000;
LUT4 lut_inst_3084 (
  .F(lut_f_3084),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_3084.INIT = 16'h8000;
LUT4 lut_inst_3085 (
  .F(lut_f_3085),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3085.INIT = 16'h8000;
LUT4 lut_inst_3086 (
  .F(lut_f_3086),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3086.INIT = 16'h8000;
LUT4 lut_inst_3087 (
  .F(lut_f_3087),
  .I0(lut_f_3084),
  .I1(lut_f_3085),
  .I2(lut_f_3086),
  .I3(gw_vcc)
);
defparam lut_inst_3087.INIT = 16'h8000;
LUT4 lut_inst_3088 (
  .F(lut_f_3088),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_3088.INIT = 16'h8000;
LUT4 lut_inst_3089 (
  .F(lut_f_3089),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3089.INIT = 16'h8000;
LUT4 lut_inst_3090 (
  .F(lut_f_3090),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3090.INIT = 16'h8000;
LUT4 lut_inst_3091 (
  .F(lut_f_3091),
  .I0(lut_f_3088),
  .I1(lut_f_3089),
  .I2(lut_f_3090),
  .I3(gw_vcc)
);
defparam lut_inst_3091.INIT = 16'h8000;
LUT4 lut_inst_3092 (
  .F(lut_f_3092),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_3092.INIT = 16'h8000;
LUT4 lut_inst_3093 (
  .F(lut_f_3093),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3093.INIT = 16'h8000;
LUT4 lut_inst_3094 (
  .F(lut_f_3094),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3094.INIT = 16'h8000;
LUT4 lut_inst_3095 (
  .F(lut_f_3095),
  .I0(lut_f_3092),
  .I1(lut_f_3093),
  .I2(lut_f_3094),
  .I3(gw_vcc)
);
defparam lut_inst_3095.INIT = 16'h8000;
LUT4 lut_inst_3096 (
  .F(lut_f_3096),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3096.INIT = 16'h8000;
LUT4 lut_inst_3097 (
  .F(lut_f_3097),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3097.INIT = 16'h8000;
LUT4 lut_inst_3098 (
  .F(lut_f_3098),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3098.INIT = 16'h8000;
LUT4 lut_inst_3099 (
  .F(lut_f_3099),
  .I0(lut_f_3096),
  .I1(lut_f_3097),
  .I2(lut_f_3098),
  .I3(gw_vcc)
);
defparam lut_inst_3099.INIT = 16'h8000;
LUT4 lut_inst_3100 (
  .F(lut_f_3100),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3100.INIT = 16'h8000;
LUT4 lut_inst_3101 (
  .F(lut_f_3101),
  .I0(ad7_inv),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3101.INIT = 16'h8000;
LUT4 lut_inst_3102 (
  .F(lut_f_3102),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3102.INIT = 16'h8000;
LUT4 lut_inst_3103 (
  .F(lut_f_3103),
  .I0(lut_f_3100),
  .I1(lut_f_3101),
  .I2(lut_f_3102),
  .I3(gw_vcc)
);
defparam lut_inst_3103.INIT = 16'h8000;
LUT4 lut_inst_3104 (
  .F(lut_f_3104),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_3104.INIT = 16'h8000;
LUT4 lut_inst_3105 (
  .F(lut_f_3105),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3105.INIT = 16'h8000;
LUT4 lut_inst_3106 (
  .F(lut_f_3106),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3106.INIT = 16'h8000;
LUT4 lut_inst_3107 (
  .F(lut_f_3107),
  .I0(lut_f_3104),
  .I1(lut_f_3105),
  .I2(lut_f_3106),
  .I3(gw_vcc)
);
defparam lut_inst_3107.INIT = 16'h8000;
LUT4 lut_inst_3108 (
  .F(lut_f_3108),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_3108.INIT = 16'h8000;
LUT4 lut_inst_3109 (
  .F(lut_f_3109),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3109.INIT = 16'h8000;
LUT4 lut_inst_3110 (
  .F(lut_f_3110),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3110.INIT = 16'h8000;
LUT4 lut_inst_3111 (
  .F(lut_f_3111),
  .I0(lut_f_3108),
  .I1(lut_f_3109),
  .I2(lut_f_3110),
  .I3(gw_vcc)
);
defparam lut_inst_3111.INIT = 16'h8000;
LUT4 lut_inst_3112 (
  .F(lut_f_3112),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_3112.INIT = 16'h8000;
LUT4 lut_inst_3113 (
  .F(lut_f_3113),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3113.INIT = 16'h8000;
LUT4 lut_inst_3114 (
  .F(lut_f_3114),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3114.INIT = 16'h8000;
LUT4 lut_inst_3115 (
  .F(lut_f_3115),
  .I0(lut_f_3112),
  .I1(lut_f_3113),
  .I2(lut_f_3114),
  .I3(gw_vcc)
);
defparam lut_inst_3115.INIT = 16'h8000;
LUT4 lut_inst_3116 (
  .F(lut_f_3116),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_3116.INIT = 16'h8000;
LUT4 lut_inst_3117 (
  .F(lut_f_3117),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3117.INIT = 16'h8000;
LUT4 lut_inst_3118 (
  .F(lut_f_3118),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3118.INIT = 16'h8000;
LUT4 lut_inst_3119 (
  .F(lut_f_3119),
  .I0(lut_f_3116),
  .I1(lut_f_3117),
  .I2(lut_f_3118),
  .I3(gw_vcc)
);
defparam lut_inst_3119.INIT = 16'h8000;
LUT4 lut_inst_3120 (
  .F(lut_f_3120),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_3120.INIT = 16'h8000;
LUT4 lut_inst_3121 (
  .F(lut_f_3121),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3121.INIT = 16'h8000;
LUT4 lut_inst_3122 (
  .F(lut_f_3122),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3122.INIT = 16'h8000;
LUT4 lut_inst_3123 (
  .F(lut_f_3123),
  .I0(lut_f_3120),
  .I1(lut_f_3121),
  .I2(lut_f_3122),
  .I3(gw_vcc)
);
defparam lut_inst_3123.INIT = 16'h8000;
LUT4 lut_inst_3124 (
  .F(lut_f_3124),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_3124.INIT = 16'h8000;
LUT4 lut_inst_3125 (
  .F(lut_f_3125),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3125.INIT = 16'h8000;
LUT4 lut_inst_3126 (
  .F(lut_f_3126),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3126.INIT = 16'h8000;
LUT4 lut_inst_3127 (
  .F(lut_f_3127),
  .I0(lut_f_3124),
  .I1(lut_f_3125),
  .I2(lut_f_3126),
  .I3(gw_vcc)
);
defparam lut_inst_3127.INIT = 16'h8000;
LUT4 lut_inst_3128 (
  .F(lut_f_3128),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3128.INIT = 16'h8000;
LUT4 lut_inst_3129 (
  .F(lut_f_3129),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3129.INIT = 16'h8000;
LUT4 lut_inst_3130 (
  .F(lut_f_3130),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3130.INIT = 16'h8000;
LUT4 lut_inst_3131 (
  .F(lut_f_3131),
  .I0(lut_f_3128),
  .I1(lut_f_3129),
  .I2(lut_f_3130),
  .I3(gw_vcc)
);
defparam lut_inst_3131.INIT = 16'h8000;
LUT4 lut_inst_3132 (
  .F(lut_f_3132),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3132.INIT = 16'h8000;
LUT4 lut_inst_3133 (
  .F(lut_f_3133),
  .I0(ad[7]),
  .I1(ad8_inv),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3133.INIT = 16'h8000;
LUT4 lut_inst_3134 (
  .F(lut_f_3134),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3134.INIT = 16'h8000;
LUT4 lut_inst_3135 (
  .F(lut_f_3135),
  .I0(lut_f_3132),
  .I1(lut_f_3133),
  .I2(lut_f_3134),
  .I3(gw_vcc)
);
defparam lut_inst_3135.INIT = 16'h8000;
LUT4 lut_inst_3136 (
  .F(lut_f_3136),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_3136.INIT = 16'h8000;
LUT4 lut_inst_3137 (
  .F(lut_f_3137),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3137.INIT = 16'h8000;
LUT4 lut_inst_3138 (
  .F(lut_f_3138),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3138.INIT = 16'h8000;
LUT4 lut_inst_3139 (
  .F(lut_f_3139),
  .I0(lut_f_3136),
  .I1(lut_f_3137),
  .I2(lut_f_3138),
  .I3(gw_vcc)
);
defparam lut_inst_3139.INIT = 16'h8000;
LUT4 lut_inst_3140 (
  .F(lut_f_3140),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_3140.INIT = 16'h8000;
LUT4 lut_inst_3141 (
  .F(lut_f_3141),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3141.INIT = 16'h8000;
LUT4 lut_inst_3142 (
  .F(lut_f_3142),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3142.INIT = 16'h8000;
LUT4 lut_inst_3143 (
  .F(lut_f_3143),
  .I0(lut_f_3140),
  .I1(lut_f_3141),
  .I2(lut_f_3142),
  .I3(gw_vcc)
);
defparam lut_inst_3143.INIT = 16'h8000;
LUT4 lut_inst_3144 (
  .F(lut_f_3144),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_3144.INIT = 16'h8000;
LUT4 lut_inst_3145 (
  .F(lut_f_3145),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3145.INIT = 16'h8000;
LUT4 lut_inst_3146 (
  .F(lut_f_3146),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3146.INIT = 16'h8000;
LUT4 lut_inst_3147 (
  .F(lut_f_3147),
  .I0(lut_f_3144),
  .I1(lut_f_3145),
  .I2(lut_f_3146),
  .I3(gw_vcc)
);
defparam lut_inst_3147.INIT = 16'h8000;
LUT4 lut_inst_3148 (
  .F(lut_f_3148),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_3148.INIT = 16'h8000;
LUT4 lut_inst_3149 (
  .F(lut_f_3149),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3149.INIT = 16'h8000;
LUT4 lut_inst_3150 (
  .F(lut_f_3150),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3150.INIT = 16'h8000;
LUT4 lut_inst_3151 (
  .F(lut_f_3151),
  .I0(lut_f_3148),
  .I1(lut_f_3149),
  .I2(lut_f_3150),
  .I3(gw_vcc)
);
defparam lut_inst_3151.INIT = 16'h8000;
LUT4 lut_inst_3152 (
  .F(lut_f_3152),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_3152.INIT = 16'h8000;
LUT4 lut_inst_3153 (
  .F(lut_f_3153),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3153.INIT = 16'h8000;
LUT4 lut_inst_3154 (
  .F(lut_f_3154),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3154.INIT = 16'h8000;
LUT4 lut_inst_3155 (
  .F(lut_f_3155),
  .I0(lut_f_3152),
  .I1(lut_f_3153),
  .I2(lut_f_3154),
  .I3(gw_vcc)
);
defparam lut_inst_3155.INIT = 16'h8000;
LUT4 lut_inst_3156 (
  .F(lut_f_3156),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_3156.INIT = 16'h8000;
LUT4 lut_inst_3157 (
  .F(lut_f_3157),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3157.INIT = 16'h8000;
LUT4 lut_inst_3158 (
  .F(lut_f_3158),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3158.INIT = 16'h8000;
LUT4 lut_inst_3159 (
  .F(lut_f_3159),
  .I0(lut_f_3156),
  .I1(lut_f_3157),
  .I2(lut_f_3158),
  .I3(gw_vcc)
);
defparam lut_inst_3159.INIT = 16'h8000;
LUT4 lut_inst_3160 (
  .F(lut_f_3160),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3160.INIT = 16'h8000;
LUT4 lut_inst_3161 (
  .F(lut_f_3161),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3161.INIT = 16'h8000;
LUT4 lut_inst_3162 (
  .F(lut_f_3162),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3162.INIT = 16'h8000;
LUT4 lut_inst_3163 (
  .F(lut_f_3163),
  .I0(lut_f_3160),
  .I1(lut_f_3161),
  .I2(lut_f_3162),
  .I3(gw_vcc)
);
defparam lut_inst_3163.INIT = 16'h8000;
LUT4 lut_inst_3164 (
  .F(lut_f_3164),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3164.INIT = 16'h8000;
LUT4 lut_inst_3165 (
  .F(lut_f_3165),
  .I0(ad7_inv),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3165.INIT = 16'h8000;
LUT4 lut_inst_3166 (
  .F(lut_f_3166),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3166.INIT = 16'h8000;
LUT4 lut_inst_3167 (
  .F(lut_f_3167),
  .I0(lut_f_3164),
  .I1(lut_f_3165),
  .I2(lut_f_3166),
  .I3(gw_vcc)
);
defparam lut_inst_3167.INIT = 16'h8000;
LUT4 lut_inst_3168 (
  .F(lut_f_3168),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_3168.INIT = 16'h8000;
LUT4 lut_inst_3169 (
  .F(lut_f_3169),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3169.INIT = 16'h8000;
LUT4 lut_inst_3170 (
  .F(lut_f_3170),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3170.INIT = 16'h8000;
LUT4 lut_inst_3171 (
  .F(lut_f_3171),
  .I0(lut_f_3168),
  .I1(lut_f_3169),
  .I2(lut_f_3170),
  .I3(gw_vcc)
);
defparam lut_inst_3171.INIT = 16'h8000;
LUT4 lut_inst_3172 (
  .F(lut_f_3172),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad6_inv)
);
defparam lut_inst_3172.INIT = 16'h8000;
LUT4 lut_inst_3173 (
  .F(lut_f_3173),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3173.INIT = 16'h8000;
LUT4 lut_inst_3174 (
  .F(lut_f_3174),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3174.INIT = 16'h8000;
LUT4 lut_inst_3175 (
  .F(lut_f_3175),
  .I0(lut_f_3172),
  .I1(lut_f_3173),
  .I2(lut_f_3174),
  .I3(gw_vcc)
);
defparam lut_inst_3175.INIT = 16'h8000;
LUT4 lut_inst_3176 (
  .F(lut_f_3176),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_3176.INIT = 16'h8000;
LUT4 lut_inst_3177 (
  .F(lut_f_3177),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3177.INIT = 16'h8000;
LUT4 lut_inst_3178 (
  .F(lut_f_3178),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3178.INIT = 16'h8000;
LUT4 lut_inst_3179 (
  .F(lut_f_3179),
  .I0(lut_f_3176),
  .I1(lut_f_3177),
  .I2(lut_f_3178),
  .I3(gw_vcc)
);
defparam lut_inst_3179.INIT = 16'h8000;
LUT4 lut_inst_3180 (
  .F(lut_f_3180),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad6_inv)
);
defparam lut_inst_3180.INIT = 16'h8000;
LUT4 lut_inst_3181 (
  .F(lut_f_3181),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3181.INIT = 16'h8000;
LUT4 lut_inst_3182 (
  .F(lut_f_3182),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3182.INIT = 16'h8000;
LUT4 lut_inst_3183 (
  .F(lut_f_3183),
  .I0(lut_f_3180),
  .I1(lut_f_3181),
  .I2(lut_f_3182),
  .I3(gw_vcc)
);
defparam lut_inst_3183.INIT = 16'h8000;
LUT4 lut_inst_3184 (
  .F(lut_f_3184),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_3184.INIT = 16'h8000;
LUT4 lut_inst_3185 (
  .F(lut_f_3185),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3185.INIT = 16'h8000;
LUT4 lut_inst_3186 (
  .F(lut_f_3186),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3186.INIT = 16'h8000;
LUT4 lut_inst_3187 (
  .F(lut_f_3187),
  .I0(lut_f_3184),
  .I1(lut_f_3185),
  .I2(lut_f_3186),
  .I3(gw_vcc)
);
defparam lut_inst_3187.INIT = 16'h8000;
LUT4 lut_inst_3188 (
  .F(lut_f_3188),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad5_inv),
  .I3(ad[6])
);
defparam lut_inst_3188.INIT = 16'h8000;
LUT4 lut_inst_3189 (
  .F(lut_f_3189),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3189.INIT = 16'h8000;
LUT4 lut_inst_3190 (
  .F(lut_f_3190),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3190.INIT = 16'h8000;
LUT4 lut_inst_3191 (
  .F(lut_f_3191),
  .I0(lut_f_3188),
  .I1(lut_f_3189),
  .I2(lut_f_3190),
  .I3(gw_vcc)
);
defparam lut_inst_3191.INIT = 16'h8000;
LUT4 lut_inst_3192 (
  .F(lut_f_3192),
  .I0(wre),
  .I1(ad4_inv),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3192.INIT = 16'h8000;
LUT4 lut_inst_3193 (
  .F(lut_f_3193),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3193.INIT = 16'h8000;
LUT4 lut_inst_3194 (
  .F(lut_f_3194),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3194.INIT = 16'h8000;
LUT4 lut_inst_3195 (
  .F(lut_f_3195),
  .I0(lut_f_3192),
  .I1(lut_f_3193),
  .I2(lut_f_3194),
  .I3(gw_vcc)
);
defparam lut_inst_3195.INIT = 16'h8000;
LUT4 lut_inst_3196 (
  .F(lut_f_3196),
  .I0(wre),
  .I1(ad[4]),
  .I2(ad[5]),
  .I3(ad[6])
);
defparam lut_inst_3196.INIT = 16'h8000;
LUT4 lut_inst_3197 (
  .F(lut_f_3197),
  .I0(ad[7]),
  .I1(ad[8]),
  .I2(ad9_inv),
  .I3(ad10_inv)
);
defparam lut_inst_3197.INIT = 16'h8000;
LUT4 lut_inst_3198 (
  .F(lut_f_3198),
  .I0(ad11_inv),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(gw_vcc)
);
defparam lut_inst_3198.INIT = 16'h8000;
LUT4 lut_inst_3199 (
  .F(lut_f_3199),
  .I0(lut_f_3196),
  .I1(lut_f_3197),
  .I2(lut_f_3198),
  .I3(gw_vcc)
);
defparam lut_inst_3199.INIT = 16'h8000;
RAM16S4 ram16s_inst_0 (
    .DO(ram16s_inst_0_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3),
    .CLK(clk)
);

defparam ram16s_inst_0.INIT_0 = 16'h0000;
defparam ram16s_inst_0.INIT_1 = 16'h0000;
defparam ram16s_inst_0.INIT_2 = 16'h0000;
defparam ram16s_inst_0.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_1 (
    .DO(ram16s_inst_1_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_7),
    .CLK(clk)
);

defparam ram16s_inst_1.INIT_0 = 16'h0000;
defparam ram16s_inst_1.INIT_1 = 16'h0000;
defparam ram16s_inst_1.INIT_2 = 16'h0000;
defparam ram16s_inst_1.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_2 (
    .DO(ram16s_inst_2_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_11),
    .CLK(clk)
);

defparam ram16s_inst_2.INIT_0 = 16'h0000;
defparam ram16s_inst_2.INIT_1 = 16'h0000;
defparam ram16s_inst_2.INIT_2 = 16'h0000;
defparam ram16s_inst_2.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_3 (
    .DO(ram16s_inst_3_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_15),
    .CLK(clk)
);

defparam ram16s_inst_3.INIT_0 = 16'h0000;
defparam ram16s_inst_3.INIT_1 = 16'h0000;
defparam ram16s_inst_3.INIT_2 = 16'h0000;
defparam ram16s_inst_3.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_4 (
    .DO(ram16s_inst_4_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_19),
    .CLK(clk)
);

defparam ram16s_inst_4.INIT_0 = 16'h0000;
defparam ram16s_inst_4.INIT_1 = 16'h0000;
defparam ram16s_inst_4.INIT_2 = 16'h0000;
defparam ram16s_inst_4.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_5 (
    .DO(ram16s_inst_5_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_23),
    .CLK(clk)
);

defparam ram16s_inst_5.INIT_0 = 16'h0000;
defparam ram16s_inst_5.INIT_1 = 16'h0000;
defparam ram16s_inst_5.INIT_2 = 16'h0000;
defparam ram16s_inst_5.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_6 (
    .DO(ram16s_inst_6_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_27),
    .CLK(clk)
);

defparam ram16s_inst_6.INIT_0 = 16'h0000;
defparam ram16s_inst_6.INIT_1 = 16'h0000;
defparam ram16s_inst_6.INIT_2 = 16'h0000;
defparam ram16s_inst_6.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_7 (
    .DO(ram16s_inst_7_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_31),
    .CLK(clk)
);

defparam ram16s_inst_7.INIT_0 = 16'h0000;
defparam ram16s_inst_7.INIT_1 = 16'h0000;
defparam ram16s_inst_7.INIT_2 = 16'h0000;
defparam ram16s_inst_7.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_8 (
    .DO(ram16s_inst_8_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_35),
    .CLK(clk)
);

defparam ram16s_inst_8.INIT_0 = 16'h0000;
defparam ram16s_inst_8.INIT_1 = 16'h0000;
defparam ram16s_inst_8.INIT_2 = 16'h0000;
defparam ram16s_inst_8.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_9 (
    .DO(ram16s_inst_9_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_39),
    .CLK(clk)
);

defparam ram16s_inst_9.INIT_0 = 16'h0000;
defparam ram16s_inst_9.INIT_1 = 16'h0000;
defparam ram16s_inst_9.INIT_2 = 16'h0000;
defparam ram16s_inst_9.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_10 (
    .DO(ram16s_inst_10_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_43),
    .CLK(clk)
);

defparam ram16s_inst_10.INIT_0 = 16'h0000;
defparam ram16s_inst_10.INIT_1 = 16'h0000;
defparam ram16s_inst_10.INIT_2 = 16'h0000;
defparam ram16s_inst_10.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_11 (
    .DO(ram16s_inst_11_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_47),
    .CLK(clk)
);

defparam ram16s_inst_11.INIT_0 = 16'h0000;
defparam ram16s_inst_11.INIT_1 = 16'h0000;
defparam ram16s_inst_11.INIT_2 = 16'h0000;
defparam ram16s_inst_11.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_12 (
    .DO(ram16s_inst_12_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_51),
    .CLK(clk)
);

defparam ram16s_inst_12.INIT_0 = 16'h0000;
defparam ram16s_inst_12.INIT_1 = 16'h0000;
defparam ram16s_inst_12.INIT_2 = 16'h0000;
defparam ram16s_inst_12.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_13 (
    .DO(ram16s_inst_13_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_55),
    .CLK(clk)
);

defparam ram16s_inst_13.INIT_0 = 16'h0000;
defparam ram16s_inst_13.INIT_1 = 16'h0000;
defparam ram16s_inst_13.INIT_2 = 16'h0000;
defparam ram16s_inst_13.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_14 (
    .DO(ram16s_inst_14_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_59),
    .CLK(clk)
);

defparam ram16s_inst_14.INIT_0 = 16'h0000;
defparam ram16s_inst_14.INIT_1 = 16'h0000;
defparam ram16s_inst_14.INIT_2 = 16'h0000;
defparam ram16s_inst_14.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_15 (
    .DO(ram16s_inst_15_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_63),
    .CLK(clk)
);

defparam ram16s_inst_15.INIT_0 = 16'hFFF8;
defparam ram16s_inst_15.INIT_1 = 16'h0000;
defparam ram16s_inst_15.INIT_2 = 16'h0000;
defparam ram16s_inst_15.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_16 (
    .DO(ram16s_inst_16_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_67),
    .CLK(clk)
);

defparam ram16s_inst_16.INIT_0 = 16'hFFFF;
defparam ram16s_inst_16.INIT_1 = 16'h0000;
defparam ram16s_inst_16.INIT_2 = 16'h0000;
defparam ram16s_inst_16.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_17 (
    .DO(ram16s_inst_17_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_71),
    .CLK(clk)
);

defparam ram16s_inst_17.INIT_0 = 16'hFFFF;
defparam ram16s_inst_17.INIT_1 = 16'h0000;
defparam ram16s_inst_17.INIT_2 = 16'h0000;
defparam ram16s_inst_17.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_18 (
    .DO(ram16s_inst_18_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_75),
    .CLK(clk)
);

defparam ram16s_inst_18.INIT_0 = 16'hFFFF;
defparam ram16s_inst_18.INIT_1 = 16'h0000;
defparam ram16s_inst_18.INIT_2 = 16'h0000;
defparam ram16s_inst_18.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_19 (
    .DO(ram16s_inst_19_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_79),
    .CLK(clk)
);

defparam ram16s_inst_19.INIT_0 = 16'h1FFF;
defparam ram16s_inst_19.INIT_1 = 16'h0000;
defparam ram16s_inst_19.INIT_2 = 16'h0000;
defparam ram16s_inst_19.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_20 (
    .DO(ram16s_inst_20_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_83),
    .CLK(clk)
);

defparam ram16s_inst_20.INIT_0 = 16'hFFF8;
defparam ram16s_inst_20.INIT_1 = 16'h0000;
defparam ram16s_inst_20.INIT_2 = 16'h0000;
defparam ram16s_inst_20.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_21 (
    .DO(ram16s_inst_21_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_87),
    .CLK(clk)
);

defparam ram16s_inst_21.INIT_0 = 16'hFFFF;
defparam ram16s_inst_21.INIT_1 = 16'h0000;
defparam ram16s_inst_21.INIT_2 = 16'h0000;
defparam ram16s_inst_21.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_22 (
    .DO(ram16s_inst_22_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_91),
    .CLK(clk)
);

defparam ram16s_inst_22.INIT_0 = 16'hFFFF;
defparam ram16s_inst_22.INIT_1 = 16'h0000;
defparam ram16s_inst_22.INIT_2 = 16'h0000;
defparam ram16s_inst_22.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_23 (
    .DO(ram16s_inst_23_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_95),
    .CLK(clk)
);

defparam ram16s_inst_23.INIT_0 = 16'hFFFF;
defparam ram16s_inst_23.INIT_1 = 16'h0000;
defparam ram16s_inst_23.INIT_2 = 16'h0000;
defparam ram16s_inst_23.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_24 (
    .DO(ram16s_inst_24_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_99),
    .CLK(clk)
);

defparam ram16s_inst_24.INIT_0 = 16'h1FFF;
defparam ram16s_inst_24.INIT_1 = 16'h0000;
defparam ram16s_inst_24.INIT_2 = 16'h0000;
defparam ram16s_inst_24.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_25 (
    .DO(ram16s_inst_25_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_103),
    .CLK(clk)
);

defparam ram16s_inst_25.INIT_0 = 16'hFFF8;
defparam ram16s_inst_25.INIT_1 = 16'h0000;
defparam ram16s_inst_25.INIT_2 = 16'h0000;
defparam ram16s_inst_25.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_26 (
    .DO(ram16s_inst_26_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_107),
    .CLK(clk)
);

defparam ram16s_inst_26.INIT_0 = 16'hFFFF;
defparam ram16s_inst_26.INIT_1 = 16'h0000;
defparam ram16s_inst_26.INIT_2 = 16'h0000;
defparam ram16s_inst_26.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_27 (
    .DO(ram16s_inst_27_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_111),
    .CLK(clk)
);

defparam ram16s_inst_27.INIT_0 = 16'hFFFF;
defparam ram16s_inst_27.INIT_1 = 16'h0000;
defparam ram16s_inst_27.INIT_2 = 16'h0000;
defparam ram16s_inst_27.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_28 (
    .DO(ram16s_inst_28_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_115),
    .CLK(clk)
);

defparam ram16s_inst_28.INIT_0 = 16'hFFFF;
defparam ram16s_inst_28.INIT_1 = 16'h0000;
defparam ram16s_inst_28.INIT_2 = 16'h0000;
defparam ram16s_inst_28.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_29 (
    .DO(ram16s_inst_29_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_119),
    .CLK(clk)
);

defparam ram16s_inst_29.INIT_0 = 16'h1FFF;
defparam ram16s_inst_29.INIT_1 = 16'h0000;
defparam ram16s_inst_29.INIT_2 = 16'h0000;
defparam ram16s_inst_29.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_30 (
    .DO(ram16s_inst_30_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_123),
    .CLK(clk)
);

defparam ram16s_inst_30.INIT_0 = 16'hFFF8;
defparam ram16s_inst_30.INIT_1 = 16'h0000;
defparam ram16s_inst_30.INIT_2 = 16'h0000;
defparam ram16s_inst_30.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_31 (
    .DO(ram16s_inst_31_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_127),
    .CLK(clk)
);

defparam ram16s_inst_31.INIT_0 = 16'hFFFF;
defparam ram16s_inst_31.INIT_1 = 16'h0000;
defparam ram16s_inst_31.INIT_2 = 16'h0000;
defparam ram16s_inst_31.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_32 (
    .DO(ram16s_inst_32_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_131),
    .CLK(clk)
);

defparam ram16s_inst_32.INIT_0 = 16'hFFFF;
defparam ram16s_inst_32.INIT_1 = 16'h0000;
defparam ram16s_inst_32.INIT_2 = 16'h0000;
defparam ram16s_inst_32.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_33 (
    .DO(ram16s_inst_33_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_135),
    .CLK(clk)
);

defparam ram16s_inst_33.INIT_0 = 16'hFFFF;
defparam ram16s_inst_33.INIT_1 = 16'h0000;
defparam ram16s_inst_33.INIT_2 = 16'h0000;
defparam ram16s_inst_33.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_34 (
    .DO(ram16s_inst_34_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_139),
    .CLK(clk)
);

defparam ram16s_inst_34.INIT_0 = 16'h1FFF;
defparam ram16s_inst_34.INIT_1 = 16'h0000;
defparam ram16s_inst_34.INIT_2 = 16'h0000;
defparam ram16s_inst_34.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_35 (
    .DO(ram16s_inst_35_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_143),
    .CLK(clk)
);

defparam ram16s_inst_35.INIT_0 = 16'hFFF8;
defparam ram16s_inst_35.INIT_1 = 16'h0000;
defparam ram16s_inst_35.INIT_2 = 16'h0000;
defparam ram16s_inst_35.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_36 (
    .DO(ram16s_inst_36_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_147),
    .CLK(clk)
);

defparam ram16s_inst_36.INIT_0 = 16'hFFFF;
defparam ram16s_inst_36.INIT_1 = 16'h0000;
defparam ram16s_inst_36.INIT_2 = 16'h0000;
defparam ram16s_inst_36.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_37 (
    .DO(ram16s_inst_37_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_151),
    .CLK(clk)
);

defparam ram16s_inst_37.INIT_0 = 16'hFFFF;
defparam ram16s_inst_37.INIT_1 = 16'h0000;
defparam ram16s_inst_37.INIT_2 = 16'h0000;
defparam ram16s_inst_37.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_38 (
    .DO(ram16s_inst_38_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_155),
    .CLK(clk)
);

defparam ram16s_inst_38.INIT_0 = 16'hFFFF;
defparam ram16s_inst_38.INIT_1 = 16'h0000;
defparam ram16s_inst_38.INIT_2 = 16'h0000;
defparam ram16s_inst_38.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_39 (
    .DO(ram16s_inst_39_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_159),
    .CLK(clk)
);

defparam ram16s_inst_39.INIT_0 = 16'h1FFF;
defparam ram16s_inst_39.INIT_1 = 16'h0000;
defparam ram16s_inst_39.INIT_2 = 16'h0000;
defparam ram16s_inst_39.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_40 (
    .DO(ram16s_inst_40_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_163),
    .CLK(clk)
);

defparam ram16s_inst_40.INIT_0 = 16'hFFF8;
defparam ram16s_inst_40.INIT_1 = 16'h0000;
defparam ram16s_inst_40.INIT_2 = 16'h0000;
defparam ram16s_inst_40.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_41 (
    .DO(ram16s_inst_41_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_167),
    .CLK(clk)
);

defparam ram16s_inst_41.INIT_0 = 16'hFFFF;
defparam ram16s_inst_41.INIT_1 = 16'h0000;
defparam ram16s_inst_41.INIT_2 = 16'h0000;
defparam ram16s_inst_41.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_42 (
    .DO(ram16s_inst_42_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_171),
    .CLK(clk)
);

defparam ram16s_inst_42.INIT_0 = 16'hFFFF;
defparam ram16s_inst_42.INIT_1 = 16'h0000;
defparam ram16s_inst_42.INIT_2 = 16'h0000;
defparam ram16s_inst_42.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_43 (
    .DO(ram16s_inst_43_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_175),
    .CLK(clk)
);

defparam ram16s_inst_43.INIT_0 = 16'hFFFF;
defparam ram16s_inst_43.INIT_1 = 16'h0000;
defparam ram16s_inst_43.INIT_2 = 16'h0000;
defparam ram16s_inst_43.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_44 (
    .DO(ram16s_inst_44_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_179),
    .CLK(clk)
);

defparam ram16s_inst_44.INIT_0 = 16'h1FFF;
defparam ram16s_inst_44.INIT_1 = 16'h0000;
defparam ram16s_inst_44.INIT_2 = 16'h0000;
defparam ram16s_inst_44.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_45 (
    .DO(ram16s_inst_45_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_183),
    .CLK(clk)
);

defparam ram16s_inst_45.INIT_0 = 16'hFFF8;
defparam ram16s_inst_45.INIT_1 = 16'h0000;
defparam ram16s_inst_45.INIT_2 = 16'h0000;
defparam ram16s_inst_45.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_46 (
    .DO(ram16s_inst_46_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_187),
    .CLK(clk)
);

defparam ram16s_inst_46.INIT_0 = 16'h803F;
defparam ram16s_inst_46.INIT_1 = 16'h0000;
defparam ram16s_inst_46.INIT_2 = 16'h0E00;
defparam ram16s_inst_46.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_47 (
    .DO(ram16s_inst_47_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_191),
    .CLK(clk)
);

defparam ram16s_inst_47.INIT_0 = 16'h3003;
defparam ram16s_inst_47.INIT_1 = 16'h0000;
defparam ram16s_inst_47.INIT_2 = 16'h81F8;
defparam ram16s_inst_47.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_48 (
    .DO(ram16s_inst_48_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_195),
    .CLK(clk)
);

defparam ram16s_inst_48.INIT_0 = 16'hF87C;
defparam ram16s_inst_48.INIT_1 = 16'h0000;
defparam ram16s_inst_48.INIT_2 = 16'h0301;
defparam ram16s_inst_48.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_49 (
    .DO(ram16s_inst_49_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_199),
    .CLK(clk)
);

defparam ram16s_inst_49.INIT_0 = 16'h1FFF;
defparam ram16s_inst_49.INIT_1 = 16'h0000;
defparam ram16s_inst_49.INIT_2 = 16'h0000;
defparam ram16s_inst_49.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_50 (
    .DO(ram16s_inst_50_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_203),
    .CLK(clk)
);

defparam ram16s_inst_50.INIT_0 = 16'hFFF8;
defparam ram16s_inst_50.INIT_1 = 16'h0000;
defparam ram16s_inst_50.INIT_2 = 16'h0000;
defparam ram16s_inst_50.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_51 (
    .DO(ram16s_inst_51_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_207),
    .CLK(clk)
);

defparam ram16s_inst_51.INIT_0 = 16'h000F;
defparam ram16s_inst_51.INIT_1 = 16'h0000;
defparam ram16s_inst_51.INIT_2 = 16'h7FC0;
defparam ram16s_inst_51.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_52 (
    .DO(ram16s_inst_52_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_211),
    .CLK(clk)
);

defparam ram16s_inst_52.INIT_0 = 16'h2003;
defparam ram16s_inst_52.INIT_1 = 16'h0000;
defparam ram16s_inst_52.INIT_2 = 16'h8FF8;
defparam ram16s_inst_52.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_53 (
    .DO(ram16s_inst_53_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_215),
    .CLK(clk)
);

defparam ram16s_inst_53.INIT_0 = 16'hF87C;
defparam ram16s_inst_53.INIT_1 = 16'h0000;
defparam ram16s_inst_53.INIT_2 = 16'h0301;
defparam ram16s_inst_53.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_54 (
    .DO(ram16s_inst_54_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_219),
    .CLK(clk)
);

defparam ram16s_inst_54.INIT_0 = 16'h1FFF;
defparam ram16s_inst_54.INIT_1 = 16'h0000;
defparam ram16s_inst_54.INIT_2 = 16'h0000;
defparam ram16s_inst_54.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_55 (
    .DO(ram16s_inst_55_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_223),
    .CLK(clk)
);

defparam ram16s_inst_55.INIT_0 = 16'hFFF8;
defparam ram16s_inst_55.INIT_1 = 16'h0000;
defparam ram16s_inst_55.INIT_2 = 16'h0000;
defparam ram16s_inst_55.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_56 (
    .DO(ram16s_inst_56_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_227),
    .CLK(clk)
);

defparam ram16s_inst_56.INIT_0 = 16'h040F;
defparam ram16s_inst_56.INIT_1 = 16'h0000;
defparam ram16s_inst_56.INIT_2 = 16'h40E0;
defparam ram16s_inst_56.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_57 (
    .DO(ram16s_inst_57_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_231),
    .CLK(clk)
);

defparam ram16s_inst_57.INIT_0 = 16'h20C3;
defparam ram16s_inst_57.INIT_1 = 16'h0000;
defparam ram16s_inst_57.INIT_2 = 16'h8C18;
defparam ram16s_inst_57.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_58 (
    .DO(ram16s_inst_58_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_235),
    .CLK(clk)
);

defparam ram16s_inst_58.INIT_0 = 16'hF87C;
defparam ram16s_inst_58.INIT_1 = 16'h0000;
defparam ram16s_inst_58.INIT_2 = 16'h0301;
defparam ram16s_inst_58.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_59 (
    .DO(ram16s_inst_59_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_239),
    .CLK(clk)
);

defparam ram16s_inst_59.INIT_0 = 16'h1FFF;
defparam ram16s_inst_59.INIT_1 = 16'h0000;
defparam ram16s_inst_59.INIT_2 = 16'h0000;
defparam ram16s_inst_59.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_60 (
    .DO(ram16s_inst_60_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_243),
    .CLK(clk)
);

defparam ram16s_inst_60.INIT_0 = 16'hFFF8;
defparam ram16s_inst_60.INIT_1 = 16'h0000;
defparam ram16s_inst_60.INIT_2 = 16'h0000;
defparam ram16s_inst_60.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_61 (
    .DO(ram16s_inst_61_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_247),
    .CLK(clk)
);

defparam ram16s_inst_61.INIT_0 = 16'h3F07;
defparam ram16s_inst_61.INIT_1 = 16'h0000;
defparam ram16s_inst_61.INIT_2 = 16'h0070;
defparam ram16s_inst_61.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_62 (
    .DO(ram16s_inst_62_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_251),
    .CLK(clk)
);

defparam ram16s_inst_62.INIT_0 = 16'h21C3;
defparam ram16s_inst_62.INIT_1 = 16'h0000;
defparam ram16s_inst_62.INIT_2 = 16'h9C18;
defparam ram16s_inst_62.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_63 (
    .DO(ram16s_inst_63_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_255),
    .CLK(clk)
);

defparam ram16s_inst_63.INIT_0 = 16'hF87C;
defparam ram16s_inst_63.INIT_1 = 16'h0000;
defparam ram16s_inst_63.INIT_2 = 16'h0301;
defparam ram16s_inst_63.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_64 (
    .DO(ram16s_inst_64_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_259),
    .CLK(clk)
);

defparam ram16s_inst_64.INIT_0 = 16'h1FFF;
defparam ram16s_inst_64.INIT_1 = 16'h0000;
defparam ram16s_inst_64.INIT_2 = 16'h0000;
defparam ram16s_inst_64.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_65 (
    .DO(ram16s_inst_65_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_263),
    .CLK(clk)
);

defparam ram16s_inst_65.INIT_0 = 16'hFFF8;
defparam ram16s_inst_65.INIT_1 = 16'h0000;
defparam ram16s_inst_65.INIT_2 = 16'h0000;
defparam ram16s_inst_65.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_66 (
    .DO(ram16s_inst_66_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_267),
    .CLK(clk)
);

defparam ram16s_inst_66.INIT_0 = 16'hFF87;
defparam ram16s_inst_66.INIT_1 = 16'h0000;
defparam ram16s_inst_66.INIT_2 = 16'h0030;
defparam ram16s_inst_66.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_67 (
    .DO(ram16s_inst_67_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_271),
    .CLK(clk)
);

defparam ram16s_inst_67.INIT_0 = 16'h21C3;
defparam ram16s_inst_67.INIT_1 = 16'h0000;
defparam ram16s_inst_67.INIT_2 = 16'h9C18;
defparam ram16s_inst_67.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_68 (
    .DO(ram16s_inst_68_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_275),
    .CLK(clk)
);

defparam ram16s_inst_68.INIT_0 = 16'hF87C;
defparam ram16s_inst_68.INIT_1 = 16'h0000;
defparam ram16s_inst_68.INIT_2 = 16'h0301;
defparam ram16s_inst_68.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_69 (
    .DO(ram16s_inst_69_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_279),
    .CLK(clk)
);

defparam ram16s_inst_69.INIT_0 = 16'h1FFF;
defparam ram16s_inst_69.INIT_1 = 16'h0000;
defparam ram16s_inst_69.INIT_2 = 16'h0000;
defparam ram16s_inst_69.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_70 (
    .DO(ram16s_inst_70_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_283),
    .CLK(clk)
);

defparam ram16s_inst_70.INIT_0 = 16'hFFF8;
defparam ram16s_inst_70.INIT_1 = 16'h0000;
defparam ram16s_inst_70.INIT_2 = 16'h0000;
defparam ram16s_inst_70.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_71 (
    .DO(ram16s_inst_71_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_287),
    .CLK(clk)
);

defparam ram16s_inst_71.INIT_0 = 16'hFF83;
defparam ram16s_inst_71.INIT_1 = 16'h0000;
defparam ram16s_inst_71.INIT_2 = 16'h0038;
defparam ram16s_inst_71.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_72 (
    .DO(ram16s_inst_72_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_291),
    .CLK(clk)
);

defparam ram16s_inst_72.INIT_0 = 16'h21C3;
defparam ram16s_inst_72.INIT_1 = 16'h0000;
defparam ram16s_inst_72.INIT_2 = 16'h8C18;
defparam ram16s_inst_72.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_73 (
    .DO(ram16s_inst_73_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_295),
    .CLK(clk)
);

defparam ram16s_inst_73.INIT_0 = 16'hF87C;
defparam ram16s_inst_73.INIT_1 = 16'h0000;
defparam ram16s_inst_73.INIT_2 = 16'h0301;
defparam ram16s_inst_73.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_74 (
    .DO(ram16s_inst_74_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_299),
    .CLK(clk)
);

defparam ram16s_inst_74.INIT_0 = 16'h1FFF;
defparam ram16s_inst_74.INIT_1 = 16'h0000;
defparam ram16s_inst_74.INIT_2 = 16'h0000;
defparam ram16s_inst_74.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_75 (
    .DO(ram16s_inst_75_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_303),
    .CLK(clk)
);

defparam ram16s_inst_75.INIT_0 = 16'hFFF8;
defparam ram16s_inst_75.INIT_1 = 16'h0000;
defparam ram16s_inst_75.INIT_2 = 16'h0000;
defparam ram16s_inst_75.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_76 (
    .DO(ram16s_inst_76_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_307),
    .CLK(clk)
);

defparam ram16s_inst_76.INIT_0 = 16'hFFC3;
defparam ram16s_inst_76.INIT_1 = 16'h0000;
defparam ram16s_inst_76.INIT_2 = 16'h0038;
defparam ram16s_inst_76.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_77 (
    .DO(ram16s_inst_77_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_311),
    .CLK(clk)
);

defparam ram16s_inst_77.INIT_0 = 16'h2043;
defparam ram16s_inst_77.INIT_1 = 16'h0000;
defparam ram16s_inst_77.INIT_2 = 16'h8E18;
defparam ram16s_inst_77.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_78 (
    .DO(ram16s_inst_78_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_315),
    .CLK(clk)
);

defparam ram16s_inst_78.INIT_0 = 16'hF87C;
defparam ram16s_inst_78.INIT_1 = 16'h0000;
defparam ram16s_inst_78.INIT_2 = 16'h0301;
defparam ram16s_inst_78.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_79 (
    .DO(ram16s_inst_79_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_319),
    .CLK(clk)
);

defparam ram16s_inst_79.INIT_0 = 16'h1FFF;
defparam ram16s_inst_79.INIT_1 = 16'h0000;
defparam ram16s_inst_79.INIT_2 = 16'h0000;
defparam ram16s_inst_79.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_80 (
    .DO(ram16s_inst_80_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_323),
    .CLK(clk)
);

defparam ram16s_inst_80.INIT_0 = 16'hFFF8;
defparam ram16s_inst_80.INIT_1 = 16'h0000;
defparam ram16s_inst_80.INIT_2 = 16'h0000;
defparam ram16s_inst_80.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_81 (
    .DO(ram16s_inst_81_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_327),
    .CLK(clk)
);

defparam ram16s_inst_81.INIT_0 = 16'h01C3;
defparam ram16s_inst_81.INIT_1 = 16'h0000;
defparam ram16s_inst_81.INIT_2 = 16'h7C38;
defparam ram16s_inst_81.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_82 (
    .DO(ram16s_inst_82_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_331),
    .CLK(clk)
);

defparam ram16s_inst_82.INIT_0 = 16'h3003;
defparam ram16s_inst_82.INIT_1 = 16'h0000;
defparam ram16s_inst_82.INIT_2 = 16'h87F8;
defparam ram16s_inst_82.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_83 (
    .DO(ram16s_inst_83_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_335),
    .CLK(clk)
);

defparam ram16s_inst_83.INIT_0 = 16'hF87C;
defparam ram16s_inst_83.INIT_1 = 16'h0000;
defparam ram16s_inst_83.INIT_2 = 16'h0301;
defparam ram16s_inst_83.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_84 (
    .DO(ram16s_inst_84_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_339),
    .CLK(clk)
);

defparam ram16s_inst_84.INIT_0 = 16'h1FFF;
defparam ram16s_inst_84.INIT_1 = 16'h0000;
defparam ram16s_inst_84.INIT_2 = 16'h0000;
defparam ram16s_inst_84.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_85 (
    .DO(ram16s_inst_85_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_343),
    .CLK(clk)
);

defparam ram16s_inst_85.INIT_0 = 16'hFFF8;
defparam ram16s_inst_85.INIT_1 = 16'h0000;
defparam ram16s_inst_85.INIT_2 = 16'h0000;
defparam ram16s_inst_85.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_86 (
    .DO(ram16s_inst_86_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_347),
    .CLK(clk)
);

defparam ram16s_inst_86.INIT_0 = 16'h0183;
defparam ram16s_inst_86.INIT_1 = 16'h0000;
defparam ram16s_inst_86.INIT_2 = 16'h7C38;
defparam ram16s_inst_86.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_87 (
    .DO(ram16s_inst_87_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_351),
    .CLK(clk)
);

defparam ram16s_inst_87.INIT_0 = 16'h3803;
defparam ram16s_inst_87.INIT_1 = 16'h0000;
defparam ram16s_inst_87.INIT_2 = 16'h81F8;
defparam ram16s_inst_87.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_88 (
    .DO(ram16s_inst_88_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_355),
    .CLK(clk)
);

defparam ram16s_inst_88.INIT_0 = 16'hF87C;
defparam ram16s_inst_88.INIT_1 = 16'h0000;
defparam ram16s_inst_88.INIT_2 = 16'h0301;
defparam ram16s_inst_88.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_89 (
    .DO(ram16s_inst_89_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_359),
    .CLK(clk)
);

defparam ram16s_inst_89.INIT_0 = 16'h1FFF;
defparam ram16s_inst_89.INIT_1 = 16'h0000;
defparam ram16s_inst_89.INIT_2 = 16'h0000;
defparam ram16s_inst_89.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_90 (
    .DO(ram16s_inst_90_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_363),
    .CLK(clk)
);

defparam ram16s_inst_90.INIT_0 = 16'hFFF8;
defparam ram16s_inst_90.INIT_1 = 16'h0000;
defparam ram16s_inst_90.INIT_2 = 16'h0000;
defparam ram16s_inst_90.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_91 (
    .DO(ram16s_inst_91_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_367),
    .CLK(clk)
);

defparam ram16s_inst_91.INIT_0 = 16'h0F87;
defparam ram16s_inst_91.INIT_1 = 16'h0000;
defparam ram16s_inst_91.INIT_2 = 16'h6030;
defparam ram16s_inst_91.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_92 (
    .DO(ram16s_inst_92_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_371),
    .CLK(clk)
);

defparam ram16s_inst_92.INIT_0 = 16'h3FC3;
defparam ram16s_inst_92.INIT_1 = 16'h0000;
defparam ram16s_inst_92.INIT_2 = 16'h8018;
defparam ram16s_inst_92.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_93 (
    .DO(ram16s_inst_93_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_375),
    .CLK(clk)
);

defparam ram16s_inst_93.INIT_0 = 16'hF87C;
defparam ram16s_inst_93.INIT_1 = 16'h0000;
defparam ram16s_inst_93.INIT_2 = 16'h0301;
defparam ram16s_inst_93.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_94 (
    .DO(ram16s_inst_94_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_379),
    .CLK(clk)
);

defparam ram16s_inst_94.INIT_0 = 16'h1FFF;
defparam ram16s_inst_94.INIT_1 = 16'h0000;
defparam ram16s_inst_94.INIT_2 = 16'h0000;
defparam ram16s_inst_94.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_95 (
    .DO(ram16s_inst_95_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_383),
    .CLK(clk)
);

defparam ram16s_inst_95.INIT_0 = 16'hFFF8;
defparam ram16s_inst_95.INIT_1 = 16'h0000;
defparam ram16s_inst_95.INIT_2 = 16'h0000;
defparam ram16s_inst_95.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_96 (
    .DO(ram16s_inst_96_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_387),
    .CLK(clk)
);

defparam ram16s_inst_96.INIT_0 = 16'h0F07;
defparam ram16s_inst_96.INIT_1 = 16'h0000;
defparam ram16s_inst_96.INIT_2 = 16'h6070;
defparam ram16s_inst_96.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_97 (
    .DO(ram16s_inst_97_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_391),
    .CLK(clk)
);

defparam ram16s_inst_97.INIT_0 = 16'h7FC3;
defparam ram16s_inst_97.INIT_1 = 16'h0000;
defparam ram16s_inst_97.INIT_2 = 16'h8018;
defparam ram16s_inst_97.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_98 (
    .DO(ram16s_inst_98_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_395),
    .CLK(clk)
);

defparam ram16s_inst_98.INIT_0 = 16'hF878;
defparam ram16s_inst_98.INIT_1 = 16'h0000;
defparam ram16s_inst_98.INIT_2 = 16'h0303;
defparam ram16s_inst_98.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_99 (
    .DO(ram16s_inst_99_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_399),
    .CLK(clk)
);

defparam ram16s_inst_99.INIT_0 = 16'h1FFF;
defparam ram16s_inst_99.INIT_1 = 16'h0000;
defparam ram16s_inst_99.INIT_2 = 16'h0000;
defparam ram16s_inst_99.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_100 (
    .DO(ram16s_inst_100_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_403),
    .CLK(clk)
);

defparam ram16s_inst_100.INIT_0 = 16'hFFF8;
defparam ram16s_inst_100.INIT_1 = 16'h0000;
defparam ram16s_inst_100.INIT_2 = 16'h0000;
defparam ram16s_inst_100.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_101 (
    .DO(ram16s_inst_101_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_407),
    .CLK(clk)
);

defparam ram16s_inst_101.INIT_0 = 16'h0C07;
defparam ram16s_inst_101.INIT_1 = 16'h0000;
defparam ram16s_inst_101.INIT_2 = 16'h60E0;
defparam ram16s_inst_101.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_102 (
    .DO(ram16s_inst_102_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_411),
    .CLK(clk)
);

defparam ram16s_inst_102.INIT_0 = 16'h7FC3;
defparam ram16s_inst_102.INIT_1 = 16'h0000;
defparam ram16s_inst_102.INIT_2 = 16'h0018;
defparam ram16s_inst_102.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_103 (
    .DO(ram16s_inst_103_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_415),
    .CLK(clk)
);

defparam ram16s_inst_103.INIT_0 = 16'hF810;
defparam ram16s_inst_103.INIT_1 = 16'h0000;
defparam ram16s_inst_103.INIT_2 = 16'h0383;
defparam ram16s_inst_103.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_104 (
    .DO(ram16s_inst_104_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_419),
    .CLK(clk)
);

defparam ram16s_inst_104.INIT_0 = 16'h1FFF;
defparam ram16s_inst_104.INIT_1 = 16'h0000;
defparam ram16s_inst_104.INIT_2 = 16'h0000;
defparam ram16s_inst_104.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_105 (
    .DO(ram16s_inst_105_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_423),
    .CLK(clk)
);

defparam ram16s_inst_105.INIT_0 = 16'hFFF8;
defparam ram16s_inst_105.INIT_1 = 16'h0000;
defparam ram16s_inst_105.INIT_2 = 16'h0000;
defparam ram16s_inst_105.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_106 (
    .DO(ram16s_inst_106_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_427),
    .CLK(clk)
);

defparam ram16s_inst_106.INIT_0 = 16'h000F;
defparam ram16s_inst_106.INIT_1 = 16'h0000;
defparam ram16s_inst_106.INIT_2 = 16'h7FC0;
defparam ram16s_inst_106.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_107 (
    .DO(ram16s_inst_107_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_431),
    .CLK(clk)
);

defparam ram16s_inst_107.INIT_0 = 16'h7FC3;
defparam ram16s_inst_107.INIT_1 = 16'h0000;
defparam ram16s_inst_107.INIT_2 = 16'h0018;
defparam ram16s_inst_107.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_108 (
    .DO(ram16s_inst_108_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_435),
    .CLK(clk)
);

defparam ram16s_inst_108.INIT_0 = 16'hFC00;
defparam ram16s_inst_108.INIT_1 = 16'h0000;
defparam ram16s_inst_108.INIT_2 = 16'h01FE;
defparam ram16s_inst_108.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_109 (
    .DO(ram16s_inst_109_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_439),
    .CLK(clk)
);

defparam ram16s_inst_109.INIT_0 = 16'h1FFF;
defparam ram16s_inst_109.INIT_1 = 16'h0000;
defparam ram16s_inst_109.INIT_2 = 16'h0000;
defparam ram16s_inst_109.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_110 (
    .DO(ram16s_inst_110_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_443),
    .CLK(clk)
);

defparam ram16s_inst_110.INIT_0 = 16'hFFF8;
defparam ram16s_inst_110.INIT_1 = 16'h0000;
defparam ram16s_inst_110.INIT_2 = 16'h0000;
defparam ram16s_inst_110.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_111 (
    .DO(ram16s_inst_111_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_447),
    .CLK(clk)
);

defparam ram16s_inst_111.INIT_0 = 16'h803F;
defparam ram16s_inst_111.INIT_1 = 16'h0000;
defparam ram16s_inst_111.INIT_2 = 16'h0E00;
defparam ram16s_inst_111.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_112 (
    .DO(ram16s_inst_112_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_451),
    .CLK(clk)
);

defparam ram16s_inst_112.INIT_0 = 16'hFFC3;
defparam ram16s_inst_112.INIT_1 = 16'h0000;
defparam ram16s_inst_112.INIT_2 = 16'h0018;
defparam ram16s_inst_112.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_113 (
    .DO(ram16s_inst_113_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_455),
    .CLK(clk)
);

defparam ram16s_inst_113.INIT_0 = 16'hFE01;
defparam ram16s_inst_113.INIT_1 = 16'h0000;
defparam ram16s_inst_113.INIT_2 = 16'h0038;
defparam ram16s_inst_113.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_114 (
    .DO(ram16s_inst_114_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_459),
    .CLK(clk)
);

defparam ram16s_inst_114.INIT_0 = 16'h1FFF;
defparam ram16s_inst_114.INIT_1 = 16'h0000;
defparam ram16s_inst_114.INIT_2 = 16'h0000;
defparam ram16s_inst_114.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_115 (
    .DO(ram16s_inst_115_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_463),
    .CLK(clk)
);

defparam ram16s_inst_115.INIT_0 = 16'hFFF8;
defparam ram16s_inst_115.INIT_1 = 16'h0000;
defparam ram16s_inst_115.INIT_2 = 16'h0000;
defparam ram16s_inst_115.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_116 (
    .DO(ram16s_inst_116_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_467),
    .CLK(clk)
);

defparam ram16s_inst_116.INIT_0 = 16'hFFFF;
defparam ram16s_inst_116.INIT_1 = 16'h0000;
defparam ram16s_inst_116.INIT_2 = 16'h0000;
defparam ram16s_inst_116.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_117 (
    .DO(ram16s_inst_117_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_471),
    .CLK(clk)
);

defparam ram16s_inst_117.INIT_0 = 16'hFFFF;
defparam ram16s_inst_117.INIT_1 = 16'h0000;
defparam ram16s_inst_117.INIT_2 = 16'h0000;
defparam ram16s_inst_117.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_118 (
    .DO(ram16s_inst_118_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_475),
    .CLK(clk)
);

defparam ram16s_inst_118.INIT_0 = 16'hFFFF;
defparam ram16s_inst_118.INIT_1 = 16'h0000;
defparam ram16s_inst_118.INIT_2 = 16'h0000;
defparam ram16s_inst_118.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_119 (
    .DO(ram16s_inst_119_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_479),
    .CLK(clk)
);

defparam ram16s_inst_119.INIT_0 = 16'h1FFF;
defparam ram16s_inst_119.INIT_1 = 16'h0000;
defparam ram16s_inst_119.INIT_2 = 16'h0000;
defparam ram16s_inst_119.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_120 (
    .DO(ram16s_inst_120_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_483),
    .CLK(clk)
);

defparam ram16s_inst_120.INIT_0 = 16'hFFF8;
defparam ram16s_inst_120.INIT_1 = 16'h0000;
defparam ram16s_inst_120.INIT_2 = 16'h0000;
defparam ram16s_inst_120.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_121 (
    .DO(ram16s_inst_121_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_487),
    .CLK(clk)
);

defparam ram16s_inst_121.INIT_0 = 16'hFFFF;
defparam ram16s_inst_121.INIT_1 = 16'h0000;
defparam ram16s_inst_121.INIT_2 = 16'h0000;
defparam ram16s_inst_121.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_122 (
    .DO(ram16s_inst_122_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_491),
    .CLK(clk)
);

defparam ram16s_inst_122.INIT_0 = 16'hFFFF;
defparam ram16s_inst_122.INIT_1 = 16'h0000;
defparam ram16s_inst_122.INIT_2 = 16'h0000;
defparam ram16s_inst_122.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_123 (
    .DO(ram16s_inst_123_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_495),
    .CLK(clk)
);

defparam ram16s_inst_123.INIT_0 = 16'hFFFF;
defparam ram16s_inst_123.INIT_1 = 16'h0000;
defparam ram16s_inst_123.INIT_2 = 16'h0000;
defparam ram16s_inst_123.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_124 (
    .DO(ram16s_inst_124_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_499),
    .CLK(clk)
);

defparam ram16s_inst_124.INIT_0 = 16'h1FFF;
defparam ram16s_inst_124.INIT_1 = 16'h0000;
defparam ram16s_inst_124.INIT_2 = 16'h0000;
defparam ram16s_inst_124.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_125 (
    .DO(ram16s_inst_125_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_503),
    .CLK(clk)
);

defparam ram16s_inst_125.INIT_0 = 16'hFFF8;
defparam ram16s_inst_125.INIT_1 = 16'h0000;
defparam ram16s_inst_125.INIT_2 = 16'h0000;
defparam ram16s_inst_125.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_126 (
    .DO(ram16s_inst_126_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_507),
    .CLK(clk)
);

defparam ram16s_inst_126.INIT_0 = 16'hFFFF;
defparam ram16s_inst_126.INIT_1 = 16'h0000;
defparam ram16s_inst_126.INIT_2 = 16'h0000;
defparam ram16s_inst_126.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_127 (
    .DO(ram16s_inst_127_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_511),
    .CLK(clk)
);

defparam ram16s_inst_127.INIT_0 = 16'hFFFF;
defparam ram16s_inst_127.INIT_1 = 16'h0000;
defparam ram16s_inst_127.INIT_2 = 16'h0000;
defparam ram16s_inst_127.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_128 (
    .DO(ram16s_inst_128_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_515),
    .CLK(clk)
);

defparam ram16s_inst_128.INIT_0 = 16'hFFFF;
defparam ram16s_inst_128.INIT_1 = 16'h0000;
defparam ram16s_inst_128.INIT_2 = 16'h0000;
defparam ram16s_inst_128.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_129 (
    .DO(ram16s_inst_129_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_519),
    .CLK(clk)
);

defparam ram16s_inst_129.INIT_0 = 16'h1FFF;
defparam ram16s_inst_129.INIT_1 = 16'h0000;
defparam ram16s_inst_129.INIT_2 = 16'h0000;
defparam ram16s_inst_129.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_130 (
    .DO(ram16s_inst_130_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_523),
    .CLK(clk)
);

defparam ram16s_inst_130.INIT_0 = 16'hFFF8;
defparam ram16s_inst_130.INIT_1 = 16'h0000;
defparam ram16s_inst_130.INIT_2 = 16'h0000;
defparam ram16s_inst_130.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_131 (
    .DO(ram16s_inst_131_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_527),
    .CLK(clk)
);

defparam ram16s_inst_131.INIT_0 = 16'hFFFF;
defparam ram16s_inst_131.INIT_1 = 16'h0000;
defparam ram16s_inst_131.INIT_2 = 16'h0000;
defparam ram16s_inst_131.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_132 (
    .DO(ram16s_inst_132_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_531),
    .CLK(clk)
);

defparam ram16s_inst_132.INIT_0 = 16'hFFFF;
defparam ram16s_inst_132.INIT_1 = 16'h0000;
defparam ram16s_inst_132.INIT_2 = 16'h0000;
defparam ram16s_inst_132.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_133 (
    .DO(ram16s_inst_133_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_535),
    .CLK(clk)
);

defparam ram16s_inst_133.INIT_0 = 16'hFFFF;
defparam ram16s_inst_133.INIT_1 = 16'h0000;
defparam ram16s_inst_133.INIT_2 = 16'h0000;
defparam ram16s_inst_133.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_134 (
    .DO(ram16s_inst_134_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_539),
    .CLK(clk)
);

defparam ram16s_inst_134.INIT_0 = 16'h1FFF;
defparam ram16s_inst_134.INIT_1 = 16'h0000;
defparam ram16s_inst_134.INIT_2 = 16'h0000;
defparam ram16s_inst_134.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_135 (
    .DO(ram16s_inst_135_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_543),
    .CLK(clk)
);

defparam ram16s_inst_135.INIT_0 = 16'h0000;
defparam ram16s_inst_135.INIT_1 = 16'h0000;
defparam ram16s_inst_135.INIT_2 = 16'h0000;
defparam ram16s_inst_135.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_136 (
    .DO(ram16s_inst_136_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_547),
    .CLK(clk)
);

defparam ram16s_inst_136.INIT_0 = 16'h0000;
defparam ram16s_inst_136.INIT_1 = 16'h0000;
defparam ram16s_inst_136.INIT_2 = 16'h0000;
defparam ram16s_inst_136.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_137 (
    .DO(ram16s_inst_137_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_551),
    .CLK(clk)
);

defparam ram16s_inst_137.INIT_0 = 16'h0000;
defparam ram16s_inst_137.INIT_1 = 16'h0000;
defparam ram16s_inst_137.INIT_2 = 16'h0000;
defparam ram16s_inst_137.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_138 (
    .DO(ram16s_inst_138_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_555),
    .CLK(clk)
);

defparam ram16s_inst_138.INIT_0 = 16'h0000;
defparam ram16s_inst_138.INIT_1 = 16'h0000;
defparam ram16s_inst_138.INIT_2 = 16'h0000;
defparam ram16s_inst_138.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_139 (
    .DO(ram16s_inst_139_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_559),
    .CLK(clk)
);

defparam ram16s_inst_139.INIT_0 = 16'h0000;
defparam ram16s_inst_139.INIT_1 = 16'h0000;
defparam ram16s_inst_139.INIT_2 = 16'h0000;
defparam ram16s_inst_139.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_140 (
    .DO(ram16s_inst_140_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_563),
    .CLK(clk)
);

defparam ram16s_inst_140.INIT_0 = 16'h0000;
defparam ram16s_inst_140.INIT_1 = 16'h0000;
defparam ram16s_inst_140.INIT_2 = 16'h0000;
defparam ram16s_inst_140.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_141 (
    .DO(ram16s_inst_141_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_567),
    .CLK(clk)
);

defparam ram16s_inst_141.INIT_0 = 16'h0000;
defparam ram16s_inst_141.INIT_1 = 16'h0000;
defparam ram16s_inst_141.INIT_2 = 16'h0000;
defparam ram16s_inst_141.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_142 (
    .DO(ram16s_inst_142_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_571),
    .CLK(clk)
);

defparam ram16s_inst_142.INIT_0 = 16'h0000;
defparam ram16s_inst_142.INIT_1 = 16'h0000;
defparam ram16s_inst_142.INIT_2 = 16'h0000;
defparam ram16s_inst_142.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_143 (
    .DO(ram16s_inst_143_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_575),
    .CLK(clk)
);

defparam ram16s_inst_143.INIT_0 = 16'h0000;
defparam ram16s_inst_143.INIT_1 = 16'h0000;
defparam ram16s_inst_143.INIT_2 = 16'h0000;
defparam ram16s_inst_143.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_144 (
    .DO(ram16s_inst_144_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_579),
    .CLK(clk)
);

defparam ram16s_inst_144.INIT_0 = 16'h0000;
defparam ram16s_inst_144.INIT_1 = 16'h0000;
defparam ram16s_inst_144.INIT_2 = 16'h0000;
defparam ram16s_inst_144.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_145 (
    .DO(ram16s_inst_145_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_583),
    .CLK(clk)
);

defparam ram16s_inst_145.INIT_0 = 16'h0000;
defparam ram16s_inst_145.INIT_1 = 16'h0000;
defparam ram16s_inst_145.INIT_2 = 16'h0000;
defparam ram16s_inst_145.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_146 (
    .DO(ram16s_inst_146_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_587),
    .CLK(clk)
);

defparam ram16s_inst_146.INIT_0 = 16'h0000;
defparam ram16s_inst_146.INIT_1 = 16'h0000;
defparam ram16s_inst_146.INIT_2 = 16'h0000;
defparam ram16s_inst_146.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_147 (
    .DO(ram16s_inst_147_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_591),
    .CLK(clk)
);

defparam ram16s_inst_147.INIT_0 = 16'h0000;
defparam ram16s_inst_147.INIT_1 = 16'h0000;
defparam ram16s_inst_147.INIT_2 = 16'h0000;
defparam ram16s_inst_147.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_148 (
    .DO(ram16s_inst_148_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_595),
    .CLK(clk)
);

defparam ram16s_inst_148.INIT_0 = 16'h0000;
defparam ram16s_inst_148.INIT_1 = 16'h0000;
defparam ram16s_inst_148.INIT_2 = 16'h0000;
defparam ram16s_inst_148.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_149 (
    .DO(ram16s_inst_149_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_599),
    .CLK(clk)
);

defparam ram16s_inst_149.INIT_0 = 16'h0000;
defparam ram16s_inst_149.INIT_1 = 16'h0000;
defparam ram16s_inst_149.INIT_2 = 16'h0000;
defparam ram16s_inst_149.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_150 (
    .DO(ram16s_inst_150_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_603),
    .CLK(clk)
);

defparam ram16s_inst_150.INIT_0 = 16'h0000;
defparam ram16s_inst_150.INIT_1 = 16'h0000;
defparam ram16s_inst_150.INIT_2 = 16'h0000;
defparam ram16s_inst_150.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_151 (
    .DO(ram16s_inst_151_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_607),
    .CLK(clk)
);

defparam ram16s_inst_151.INIT_0 = 16'h0000;
defparam ram16s_inst_151.INIT_1 = 16'h0000;
defparam ram16s_inst_151.INIT_2 = 16'h0000;
defparam ram16s_inst_151.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_152 (
    .DO(ram16s_inst_152_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_611),
    .CLK(clk)
);

defparam ram16s_inst_152.INIT_0 = 16'h0000;
defparam ram16s_inst_152.INIT_1 = 16'h0000;
defparam ram16s_inst_152.INIT_2 = 16'h0000;
defparam ram16s_inst_152.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_153 (
    .DO(ram16s_inst_153_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_615),
    .CLK(clk)
);

defparam ram16s_inst_153.INIT_0 = 16'h0000;
defparam ram16s_inst_153.INIT_1 = 16'h0000;
defparam ram16s_inst_153.INIT_2 = 16'h0000;
defparam ram16s_inst_153.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_154 (
    .DO(ram16s_inst_154_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_619),
    .CLK(clk)
);

defparam ram16s_inst_154.INIT_0 = 16'h0000;
defparam ram16s_inst_154.INIT_1 = 16'h0000;
defparam ram16s_inst_154.INIT_2 = 16'h0000;
defparam ram16s_inst_154.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_155 (
    .DO(ram16s_inst_155_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_623),
    .CLK(clk)
);

defparam ram16s_inst_155.INIT_0 = 16'h0000;
defparam ram16s_inst_155.INIT_1 = 16'h0000;
defparam ram16s_inst_155.INIT_2 = 16'h0000;
defparam ram16s_inst_155.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_156 (
    .DO(ram16s_inst_156_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_627),
    .CLK(clk)
);

defparam ram16s_inst_156.INIT_0 = 16'h0000;
defparam ram16s_inst_156.INIT_1 = 16'h0000;
defparam ram16s_inst_156.INIT_2 = 16'h0000;
defparam ram16s_inst_156.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_157 (
    .DO(ram16s_inst_157_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_631),
    .CLK(clk)
);

defparam ram16s_inst_157.INIT_0 = 16'h0000;
defparam ram16s_inst_157.INIT_1 = 16'h0000;
defparam ram16s_inst_157.INIT_2 = 16'h0000;
defparam ram16s_inst_157.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_158 (
    .DO(ram16s_inst_158_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_635),
    .CLK(clk)
);

defparam ram16s_inst_158.INIT_0 = 16'h0000;
defparam ram16s_inst_158.INIT_1 = 16'h0000;
defparam ram16s_inst_158.INIT_2 = 16'h0000;
defparam ram16s_inst_158.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_159 (
    .DO(ram16s_inst_159_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_639),
    .CLK(clk)
);

defparam ram16s_inst_159.INIT_0 = 16'h0000;
defparam ram16s_inst_159.INIT_1 = 16'h0000;
defparam ram16s_inst_159.INIT_2 = 16'h0000;
defparam ram16s_inst_159.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_160 (
    .DO(ram16s_inst_160_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_643),
    .CLK(clk)
);

defparam ram16s_inst_160.INIT_0 = 16'h0000;
defparam ram16s_inst_160.INIT_1 = 16'h0000;
defparam ram16s_inst_160.INIT_2 = 16'h0000;
defparam ram16s_inst_160.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_161 (
    .DO(ram16s_inst_161_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_647),
    .CLK(clk)
);

defparam ram16s_inst_161.INIT_0 = 16'h0000;
defparam ram16s_inst_161.INIT_1 = 16'h0000;
defparam ram16s_inst_161.INIT_2 = 16'h0000;
defparam ram16s_inst_161.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_162 (
    .DO(ram16s_inst_162_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_651),
    .CLK(clk)
);

defparam ram16s_inst_162.INIT_0 = 16'h0000;
defparam ram16s_inst_162.INIT_1 = 16'h0000;
defparam ram16s_inst_162.INIT_2 = 16'h0000;
defparam ram16s_inst_162.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_163 (
    .DO(ram16s_inst_163_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_655),
    .CLK(clk)
);

defparam ram16s_inst_163.INIT_0 = 16'h0000;
defparam ram16s_inst_163.INIT_1 = 16'h0000;
defparam ram16s_inst_163.INIT_2 = 16'h0000;
defparam ram16s_inst_163.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_164 (
    .DO(ram16s_inst_164_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_659),
    .CLK(clk)
);

defparam ram16s_inst_164.INIT_0 = 16'h0000;
defparam ram16s_inst_164.INIT_1 = 16'h0000;
defparam ram16s_inst_164.INIT_2 = 16'h0000;
defparam ram16s_inst_164.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_165 (
    .DO(ram16s_inst_165_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_663),
    .CLK(clk)
);

defparam ram16s_inst_165.INIT_0 = 16'h0000;
defparam ram16s_inst_165.INIT_1 = 16'h0000;
defparam ram16s_inst_165.INIT_2 = 16'h0000;
defparam ram16s_inst_165.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_166 (
    .DO(ram16s_inst_166_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_667),
    .CLK(clk)
);

defparam ram16s_inst_166.INIT_0 = 16'h0000;
defparam ram16s_inst_166.INIT_1 = 16'h0000;
defparam ram16s_inst_166.INIT_2 = 16'h0000;
defparam ram16s_inst_166.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_167 (
    .DO(ram16s_inst_167_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_671),
    .CLK(clk)
);

defparam ram16s_inst_167.INIT_0 = 16'h0000;
defparam ram16s_inst_167.INIT_1 = 16'h0000;
defparam ram16s_inst_167.INIT_2 = 16'h0000;
defparam ram16s_inst_167.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_168 (
    .DO(ram16s_inst_168_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_675),
    .CLK(clk)
);

defparam ram16s_inst_168.INIT_0 = 16'h0000;
defparam ram16s_inst_168.INIT_1 = 16'h0000;
defparam ram16s_inst_168.INIT_2 = 16'h0000;
defparam ram16s_inst_168.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_169 (
    .DO(ram16s_inst_169_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_679),
    .CLK(clk)
);

defparam ram16s_inst_169.INIT_0 = 16'h0000;
defparam ram16s_inst_169.INIT_1 = 16'h0000;
defparam ram16s_inst_169.INIT_2 = 16'h0000;
defparam ram16s_inst_169.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_170 (
    .DO(ram16s_inst_170_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_683),
    .CLK(clk)
);

defparam ram16s_inst_170.INIT_0 = 16'h0000;
defparam ram16s_inst_170.INIT_1 = 16'h0000;
defparam ram16s_inst_170.INIT_2 = 16'h0000;
defparam ram16s_inst_170.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_171 (
    .DO(ram16s_inst_171_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_687),
    .CLK(clk)
);

defparam ram16s_inst_171.INIT_0 = 16'h0000;
defparam ram16s_inst_171.INIT_1 = 16'h0000;
defparam ram16s_inst_171.INIT_2 = 16'h0000;
defparam ram16s_inst_171.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_172 (
    .DO(ram16s_inst_172_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_691),
    .CLK(clk)
);

defparam ram16s_inst_172.INIT_0 = 16'h0000;
defparam ram16s_inst_172.INIT_1 = 16'h0000;
defparam ram16s_inst_172.INIT_2 = 16'h0000;
defparam ram16s_inst_172.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_173 (
    .DO(ram16s_inst_173_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_695),
    .CLK(clk)
);

defparam ram16s_inst_173.INIT_0 = 16'h0000;
defparam ram16s_inst_173.INIT_1 = 16'h0000;
defparam ram16s_inst_173.INIT_2 = 16'h0000;
defparam ram16s_inst_173.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_174 (
    .DO(ram16s_inst_174_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_699),
    .CLK(clk)
);

defparam ram16s_inst_174.INIT_0 = 16'h0000;
defparam ram16s_inst_174.INIT_1 = 16'h0000;
defparam ram16s_inst_174.INIT_2 = 16'h0000;
defparam ram16s_inst_174.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_175 (
    .DO(ram16s_inst_175_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_703),
    .CLK(clk)
);

defparam ram16s_inst_175.INIT_0 = 16'h0000;
defparam ram16s_inst_175.INIT_1 = 16'h0000;
defparam ram16s_inst_175.INIT_2 = 16'h0000;
defparam ram16s_inst_175.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_176 (
    .DO(ram16s_inst_176_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_707),
    .CLK(clk)
);

defparam ram16s_inst_176.INIT_0 = 16'h0000;
defparam ram16s_inst_176.INIT_1 = 16'h0000;
defparam ram16s_inst_176.INIT_2 = 16'h0000;
defparam ram16s_inst_176.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_177 (
    .DO(ram16s_inst_177_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_711),
    .CLK(clk)
);

defparam ram16s_inst_177.INIT_0 = 16'h0000;
defparam ram16s_inst_177.INIT_1 = 16'h0000;
defparam ram16s_inst_177.INIT_2 = 16'h0000;
defparam ram16s_inst_177.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_178 (
    .DO(ram16s_inst_178_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_715),
    .CLK(clk)
);

defparam ram16s_inst_178.INIT_0 = 16'h0000;
defparam ram16s_inst_178.INIT_1 = 16'h0000;
defparam ram16s_inst_178.INIT_2 = 16'h0000;
defparam ram16s_inst_178.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_179 (
    .DO(ram16s_inst_179_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_719),
    .CLK(clk)
);

defparam ram16s_inst_179.INIT_0 = 16'h0000;
defparam ram16s_inst_179.INIT_1 = 16'h0000;
defparam ram16s_inst_179.INIT_2 = 16'h0000;
defparam ram16s_inst_179.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_180 (
    .DO(ram16s_inst_180_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_723),
    .CLK(clk)
);

defparam ram16s_inst_180.INIT_0 = 16'h0000;
defparam ram16s_inst_180.INIT_1 = 16'h0000;
defparam ram16s_inst_180.INIT_2 = 16'h0000;
defparam ram16s_inst_180.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_181 (
    .DO(ram16s_inst_181_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_727),
    .CLK(clk)
);

defparam ram16s_inst_181.INIT_0 = 16'h0000;
defparam ram16s_inst_181.INIT_1 = 16'h0000;
defparam ram16s_inst_181.INIT_2 = 16'h0000;
defparam ram16s_inst_181.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_182 (
    .DO(ram16s_inst_182_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_731),
    .CLK(clk)
);

defparam ram16s_inst_182.INIT_0 = 16'h0000;
defparam ram16s_inst_182.INIT_1 = 16'h0000;
defparam ram16s_inst_182.INIT_2 = 16'h0000;
defparam ram16s_inst_182.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_183 (
    .DO(ram16s_inst_183_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_735),
    .CLK(clk)
);

defparam ram16s_inst_183.INIT_0 = 16'h0000;
defparam ram16s_inst_183.INIT_1 = 16'h0000;
defparam ram16s_inst_183.INIT_2 = 16'h0000;
defparam ram16s_inst_183.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_184 (
    .DO(ram16s_inst_184_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_739),
    .CLK(clk)
);

defparam ram16s_inst_184.INIT_0 = 16'h0000;
defparam ram16s_inst_184.INIT_1 = 16'h0000;
defparam ram16s_inst_184.INIT_2 = 16'h0000;
defparam ram16s_inst_184.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_185 (
    .DO(ram16s_inst_185_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_743),
    .CLK(clk)
);

defparam ram16s_inst_185.INIT_0 = 16'h0000;
defparam ram16s_inst_185.INIT_1 = 16'h0000;
defparam ram16s_inst_185.INIT_2 = 16'h0000;
defparam ram16s_inst_185.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_186 (
    .DO(ram16s_inst_186_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_747),
    .CLK(clk)
);

defparam ram16s_inst_186.INIT_0 = 16'h0000;
defparam ram16s_inst_186.INIT_1 = 16'h0000;
defparam ram16s_inst_186.INIT_2 = 16'h0000;
defparam ram16s_inst_186.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_187 (
    .DO(ram16s_inst_187_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_751),
    .CLK(clk)
);

defparam ram16s_inst_187.INIT_0 = 16'h0000;
defparam ram16s_inst_187.INIT_1 = 16'h0000;
defparam ram16s_inst_187.INIT_2 = 16'h0000;
defparam ram16s_inst_187.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_188 (
    .DO(ram16s_inst_188_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_755),
    .CLK(clk)
);

defparam ram16s_inst_188.INIT_0 = 16'h0000;
defparam ram16s_inst_188.INIT_1 = 16'h0000;
defparam ram16s_inst_188.INIT_2 = 16'h0000;
defparam ram16s_inst_188.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_189 (
    .DO(ram16s_inst_189_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_759),
    .CLK(clk)
);

defparam ram16s_inst_189.INIT_0 = 16'h0000;
defparam ram16s_inst_189.INIT_1 = 16'h0000;
defparam ram16s_inst_189.INIT_2 = 16'h0000;
defparam ram16s_inst_189.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_190 (
    .DO(ram16s_inst_190_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_763),
    .CLK(clk)
);

defparam ram16s_inst_190.INIT_0 = 16'h0000;
defparam ram16s_inst_190.INIT_1 = 16'h0000;
defparam ram16s_inst_190.INIT_2 = 16'h0000;
defparam ram16s_inst_190.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_191 (
    .DO(ram16s_inst_191_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_767),
    .CLK(clk)
);

defparam ram16s_inst_191.INIT_0 = 16'h0000;
defparam ram16s_inst_191.INIT_1 = 16'h0000;
defparam ram16s_inst_191.INIT_2 = 16'h0000;
defparam ram16s_inst_191.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_192 (
    .DO(ram16s_inst_192_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_771),
    .CLK(clk)
);

defparam ram16s_inst_192.INIT_0 = 16'h0000;
defparam ram16s_inst_192.INIT_1 = 16'h0000;
defparam ram16s_inst_192.INIT_2 = 16'h0000;
defparam ram16s_inst_192.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_193 (
    .DO(ram16s_inst_193_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_775),
    .CLK(clk)
);

defparam ram16s_inst_193.INIT_0 = 16'h0000;
defparam ram16s_inst_193.INIT_1 = 16'h0000;
defparam ram16s_inst_193.INIT_2 = 16'h0000;
defparam ram16s_inst_193.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_194 (
    .DO(ram16s_inst_194_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_779),
    .CLK(clk)
);

defparam ram16s_inst_194.INIT_0 = 16'h0000;
defparam ram16s_inst_194.INIT_1 = 16'h0000;
defparam ram16s_inst_194.INIT_2 = 16'h0000;
defparam ram16s_inst_194.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_195 (
    .DO(ram16s_inst_195_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_783),
    .CLK(clk)
);

defparam ram16s_inst_195.INIT_0 = 16'h0000;
defparam ram16s_inst_195.INIT_1 = 16'h0000;
defparam ram16s_inst_195.INIT_2 = 16'h0000;
defparam ram16s_inst_195.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_196 (
    .DO(ram16s_inst_196_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_787),
    .CLK(clk)
);

defparam ram16s_inst_196.INIT_0 = 16'h0000;
defparam ram16s_inst_196.INIT_1 = 16'h0000;
defparam ram16s_inst_196.INIT_2 = 16'h0000;
defparam ram16s_inst_196.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_197 (
    .DO(ram16s_inst_197_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_791),
    .CLK(clk)
);

defparam ram16s_inst_197.INIT_0 = 16'h0000;
defparam ram16s_inst_197.INIT_1 = 16'h0000;
defparam ram16s_inst_197.INIT_2 = 16'h0000;
defparam ram16s_inst_197.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_198 (
    .DO(ram16s_inst_198_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_795),
    .CLK(clk)
);

defparam ram16s_inst_198.INIT_0 = 16'h0000;
defparam ram16s_inst_198.INIT_1 = 16'h0000;
defparam ram16s_inst_198.INIT_2 = 16'h0000;
defparam ram16s_inst_198.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_199 (
    .DO(ram16s_inst_199_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_799),
    .CLK(clk)
);

defparam ram16s_inst_199.INIT_0 = 16'h0000;
defparam ram16s_inst_199.INIT_1 = 16'h0000;
defparam ram16s_inst_199.INIT_2 = 16'h0000;
defparam ram16s_inst_199.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_200 (
    .DO(ram16s_inst_200_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_803),
    .CLK(clk)
);

defparam ram16s_inst_200.INIT_0 = 16'h0000;
defparam ram16s_inst_200.INIT_1 = 16'h0000;
defparam ram16s_inst_200.INIT_2 = 16'h0000;
defparam ram16s_inst_200.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_201 (
    .DO(ram16s_inst_201_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_807),
    .CLK(clk)
);

defparam ram16s_inst_201.INIT_0 = 16'h0000;
defparam ram16s_inst_201.INIT_1 = 16'h0000;
defparam ram16s_inst_201.INIT_2 = 16'h0000;
defparam ram16s_inst_201.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_202 (
    .DO(ram16s_inst_202_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_811),
    .CLK(clk)
);

defparam ram16s_inst_202.INIT_0 = 16'h0000;
defparam ram16s_inst_202.INIT_1 = 16'h0000;
defparam ram16s_inst_202.INIT_2 = 16'h0000;
defparam ram16s_inst_202.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_203 (
    .DO(ram16s_inst_203_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_815),
    .CLK(clk)
);

defparam ram16s_inst_203.INIT_0 = 16'h0000;
defparam ram16s_inst_203.INIT_1 = 16'h0000;
defparam ram16s_inst_203.INIT_2 = 16'h0000;
defparam ram16s_inst_203.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_204 (
    .DO(ram16s_inst_204_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_819),
    .CLK(clk)
);

defparam ram16s_inst_204.INIT_0 = 16'h0000;
defparam ram16s_inst_204.INIT_1 = 16'h0000;
defparam ram16s_inst_204.INIT_2 = 16'h0000;
defparam ram16s_inst_204.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_205 (
    .DO(ram16s_inst_205_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_823),
    .CLK(clk)
);

defparam ram16s_inst_205.INIT_0 = 16'h0000;
defparam ram16s_inst_205.INIT_1 = 16'h0000;
defparam ram16s_inst_205.INIT_2 = 16'h0000;
defparam ram16s_inst_205.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_206 (
    .DO(ram16s_inst_206_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_827),
    .CLK(clk)
);

defparam ram16s_inst_206.INIT_0 = 16'h0000;
defparam ram16s_inst_206.INIT_1 = 16'h0000;
defparam ram16s_inst_206.INIT_2 = 16'h0000;
defparam ram16s_inst_206.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_207 (
    .DO(ram16s_inst_207_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_831),
    .CLK(clk)
);

defparam ram16s_inst_207.INIT_0 = 16'h0000;
defparam ram16s_inst_207.INIT_1 = 16'h0000;
defparam ram16s_inst_207.INIT_2 = 16'h0000;
defparam ram16s_inst_207.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_208 (
    .DO(ram16s_inst_208_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_835),
    .CLK(clk)
);

defparam ram16s_inst_208.INIT_0 = 16'h0000;
defparam ram16s_inst_208.INIT_1 = 16'h0000;
defparam ram16s_inst_208.INIT_2 = 16'h0000;
defparam ram16s_inst_208.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_209 (
    .DO(ram16s_inst_209_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_839),
    .CLK(clk)
);

defparam ram16s_inst_209.INIT_0 = 16'h0000;
defparam ram16s_inst_209.INIT_1 = 16'h0000;
defparam ram16s_inst_209.INIT_2 = 16'h0000;
defparam ram16s_inst_209.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_210 (
    .DO(ram16s_inst_210_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_843),
    .CLK(clk)
);

defparam ram16s_inst_210.INIT_0 = 16'h0000;
defparam ram16s_inst_210.INIT_1 = 16'h0000;
defparam ram16s_inst_210.INIT_2 = 16'h0000;
defparam ram16s_inst_210.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_211 (
    .DO(ram16s_inst_211_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_847),
    .CLK(clk)
);

defparam ram16s_inst_211.INIT_0 = 16'h0000;
defparam ram16s_inst_211.INIT_1 = 16'h0000;
defparam ram16s_inst_211.INIT_2 = 16'h0000;
defparam ram16s_inst_211.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_212 (
    .DO(ram16s_inst_212_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_851),
    .CLK(clk)
);

defparam ram16s_inst_212.INIT_0 = 16'h0000;
defparam ram16s_inst_212.INIT_1 = 16'h0000;
defparam ram16s_inst_212.INIT_2 = 16'h0000;
defparam ram16s_inst_212.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_213 (
    .DO(ram16s_inst_213_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_855),
    .CLK(clk)
);

defparam ram16s_inst_213.INIT_0 = 16'h0000;
defparam ram16s_inst_213.INIT_1 = 16'h0000;
defparam ram16s_inst_213.INIT_2 = 16'h0000;
defparam ram16s_inst_213.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_214 (
    .DO(ram16s_inst_214_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_859),
    .CLK(clk)
);

defparam ram16s_inst_214.INIT_0 = 16'h0000;
defparam ram16s_inst_214.INIT_1 = 16'h0000;
defparam ram16s_inst_214.INIT_2 = 16'h0000;
defparam ram16s_inst_214.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_215 (
    .DO(ram16s_inst_215_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_863),
    .CLK(clk)
);

defparam ram16s_inst_215.INIT_0 = 16'h0000;
defparam ram16s_inst_215.INIT_1 = 16'h0000;
defparam ram16s_inst_215.INIT_2 = 16'h0000;
defparam ram16s_inst_215.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_216 (
    .DO(ram16s_inst_216_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_867),
    .CLK(clk)
);

defparam ram16s_inst_216.INIT_0 = 16'h0000;
defparam ram16s_inst_216.INIT_1 = 16'h0000;
defparam ram16s_inst_216.INIT_2 = 16'h0000;
defparam ram16s_inst_216.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_217 (
    .DO(ram16s_inst_217_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_871),
    .CLK(clk)
);

defparam ram16s_inst_217.INIT_0 = 16'h0000;
defparam ram16s_inst_217.INIT_1 = 16'h0000;
defparam ram16s_inst_217.INIT_2 = 16'h0000;
defparam ram16s_inst_217.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_218 (
    .DO(ram16s_inst_218_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_875),
    .CLK(clk)
);

defparam ram16s_inst_218.INIT_0 = 16'h0000;
defparam ram16s_inst_218.INIT_1 = 16'h0000;
defparam ram16s_inst_218.INIT_2 = 16'h0000;
defparam ram16s_inst_218.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_219 (
    .DO(ram16s_inst_219_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_879),
    .CLK(clk)
);

defparam ram16s_inst_219.INIT_0 = 16'h0000;
defparam ram16s_inst_219.INIT_1 = 16'h0000;
defparam ram16s_inst_219.INIT_2 = 16'h0000;
defparam ram16s_inst_219.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_220 (
    .DO(ram16s_inst_220_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_883),
    .CLK(clk)
);

defparam ram16s_inst_220.INIT_0 = 16'h0000;
defparam ram16s_inst_220.INIT_1 = 16'h0000;
defparam ram16s_inst_220.INIT_2 = 16'h0000;
defparam ram16s_inst_220.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_221 (
    .DO(ram16s_inst_221_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_887),
    .CLK(clk)
);

defparam ram16s_inst_221.INIT_0 = 16'h0000;
defparam ram16s_inst_221.INIT_1 = 16'h0000;
defparam ram16s_inst_221.INIT_2 = 16'h0000;
defparam ram16s_inst_221.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_222 (
    .DO(ram16s_inst_222_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_891),
    .CLK(clk)
);

defparam ram16s_inst_222.INIT_0 = 16'h0000;
defparam ram16s_inst_222.INIT_1 = 16'h0000;
defparam ram16s_inst_222.INIT_2 = 16'h0000;
defparam ram16s_inst_222.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_223 (
    .DO(ram16s_inst_223_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_895),
    .CLK(clk)
);

defparam ram16s_inst_223.INIT_0 = 16'h0000;
defparam ram16s_inst_223.INIT_1 = 16'h0000;
defparam ram16s_inst_223.INIT_2 = 16'h0000;
defparam ram16s_inst_223.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_224 (
    .DO(ram16s_inst_224_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_899),
    .CLK(clk)
);

defparam ram16s_inst_224.INIT_0 = 16'h0000;
defparam ram16s_inst_224.INIT_1 = 16'h0000;
defparam ram16s_inst_224.INIT_2 = 16'h0000;
defparam ram16s_inst_224.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_225 (
    .DO(ram16s_inst_225_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_903),
    .CLK(clk)
);

defparam ram16s_inst_225.INIT_0 = 16'h0000;
defparam ram16s_inst_225.INIT_1 = 16'h0000;
defparam ram16s_inst_225.INIT_2 = 16'h0000;
defparam ram16s_inst_225.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_226 (
    .DO(ram16s_inst_226_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_907),
    .CLK(clk)
);

defparam ram16s_inst_226.INIT_0 = 16'h0000;
defparam ram16s_inst_226.INIT_1 = 16'h0000;
defparam ram16s_inst_226.INIT_2 = 16'h0000;
defparam ram16s_inst_226.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_227 (
    .DO(ram16s_inst_227_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_911),
    .CLK(clk)
);

defparam ram16s_inst_227.INIT_0 = 16'h0000;
defparam ram16s_inst_227.INIT_1 = 16'h0000;
defparam ram16s_inst_227.INIT_2 = 16'h0000;
defparam ram16s_inst_227.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_228 (
    .DO(ram16s_inst_228_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_915),
    .CLK(clk)
);

defparam ram16s_inst_228.INIT_0 = 16'h0000;
defparam ram16s_inst_228.INIT_1 = 16'h0000;
defparam ram16s_inst_228.INIT_2 = 16'h0000;
defparam ram16s_inst_228.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_229 (
    .DO(ram16s_inst_229_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_919),
    .CLK(clk)
);

defparam ram16s_inst_229.INIT_0 = 16'h0000;
defparam ram16s_inst_229.INIT_1 = 16'h0000;
defparam ram16s_inst_229.INIT_2 = 16'h0000;
defparam ram16s_inst_229.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_230 (
    .DO(ram16s_inst_230_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_923),
    .CLK(clk)
);

defparam ram16s_inst_230.INIT_0 = 16'h0000;
defparam ram16s_inst_230.INIT_1 = 16'h0000;
defparam ram16s_inst_230.INIT_2 = 16'h0000;
defparam ram16s_inst_230.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_231 (
    .DO(ram16s_inst_231_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_927),
    .CLK(clk)
);

defparam ram16s_inst_231.INIT_0 = 16'h0000;
defparam ram16s_inst_231.INIT_1 = 16'h0000;
defparam ram16s_inst_231.INIT_2 = 16'h0000;
defparam ram16s_inst_231.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_232 (
    .DO(ram16s_inst_232_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_931),
    .CLK(clk)
);

defparam ram16s_inst_232.INIT_0 = 16'h0000;
defparam ram16s_inst_232.INIT_1 = 16'h0000;
defparam ram16s_inst_232.INIT_2 = 16'h0000;
defparam ram16s_inst_232.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_233 (
    .DO(ram16s_inst_233_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_935),
    .CLK(clk)
);

defparam ram16s_inst_233.INIT_0 = 16'h0000;
defparam ram16s_inst_233.INIT_1 = 16'h0000;
defparam ram16s_inst_233.INIT_2 = 16'h0000;
defparam ram16s_inst_233.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_234 (
    .DO(ram16s_inst_234_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_939),
    .CLK(clk)
);

defparam ram16s_inst_234.INIT_0 = 16'h0000;
defparam ram16s_inst_234.INIT_1 = 16'h0000;
defparam ram16s_inst_234.INIT_2 = 16'h0000;
defparam ram16s_inst_234.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_235 (
    .DO(ram16s_inst_235_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_943),
    .CLK(clk)
);

defparam ram16s_inst_235.INIT_0 = 16'hC000;
defparam ram16s_inst_235.INIT_1 = 16'h0000;
defparam ram16s_inst_235.INIT_2 = 16'h0000;
defparam ram16s_inst_235.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_236 (
    .DO(ram16s_inst_236_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_947),
    .CLK(clk)
);

defparam ram16s_inst_236.INIT_0 = 16'h0001;
defparam ram16s_inst_236.INIT_1 = 16'h0000;
defparam ram16s_inst_236.INIT_2 = 16'h0000;
defparam ram16s_inst_236.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_237 (
    .DO(ram16s_inst_237_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_951),
    .CLK(clk)
);

defparam ram16s_inst_237.INIT_0 = 16'h0000;
defparam ram16s_inst_237.INIT_1 = 16'h0000;
defparam ram16s_inst_237.INIT_2 = 16'h0000;
defparam ram16s_inst_237.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_238 (
    .DO(ram16s_inst_238_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_955),
    .CLK(clk)
);

defparam ram16s_inst_238.INIT_0 = 16'h0000;
defparam ram16s_inst_238.INIT_1 = 16'h0000;
defparam ram16s_inst_238.INIT_2 = 16'h0000;
defparam ram16s_inst_238.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_239 (
    .DO(ram16s_inst_239_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_959),
    .CLK(clk)
);

defparam ram16s_inst_239.INIT_0 = 16'h0000;
defparam ram16s_inst_239.INIT_1 = 16'h0000;
defparam ram16s_inst_239.INIT_2 = 16'h0000;
defparam ram16s_inst_239.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_240 (
    .DO(ram16s_inst_240_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_963),
    .CLK(clk)
);

defparam ram16s_inst_240.INIT_0 = 16'hF000;
defparam ram16s_inst_240.INIT_1 = 16'h0000;
defparam ram16s_inst_240.INIT_2 = 16'h0000;
defparam ram16s_inst_240.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_241 (
    .DO(ram16s_inst_241_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_967),
    .CLK(clk)
);

defparam ram16s_inst_241.INIT_0 = 16'h0007;
defparam ram16s_inst_241.INIT_1 = 16'h0000;
defparam ram16s_inst_241.INIT_2 = 16'h0000;
defparam ram16s_inst_241.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_242 (
    .DO(ram16s_inst_242_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_971),
    .CLK(clk)
);

defparam ram16s_inst_242.INIT_0 = 16'h0000;
defparam ram16s_inst_242.INIT_1 = 16'h0000;
defparam ram16s_inst_242.INIT_2 = 16'h0000;
defparam ram16s_inst_242.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_243 (
    .DO(ram16s_inst_243_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_975),
    .CLK(clk)
);

defparam ram16s_inst_243.INIT_0 = 16'h0000;
defparam ram16s_inst_243.INIT_1 = 16'h0000;
defparam ram16s_inst_243.INIT_2 = 16'h0000;
defparam ram16s_inst_243.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_244 (
    .DO(ram16s_inst_244_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_979),
    .CLK(clk)
);

defparam ram16s_inst_244.INIT_0 = 16'h0000;
defparam ram16s_inst_244.INIT_1 = 16'h0000;
defparam ram16s_inst_244.INIT_2 = 16'h0000;
defparam ram16s_inst_244.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_245 (
    .DO(ram16s_inst_245_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_983),
    .CLK(clk)
);

defparam ram16s_inst_245.INIT_0 = 16'h1800;
defparam ram16s_inst_245.INIT_1 = 16'h0000;
defparam ram16s_inst_245.INIT_2 = 16'h0000;
defparam ram16s_inst_245.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_246 (
    .DO(ram16s_inst_246_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_987),
    .CLK(clk)
);

defparam ram16s_inst_246.INIT_0 = 16'h0004;
defparam ram16s_inst_246.INIT_1 = 16'h0000;
defparam ram16s_inst_246.INIT_2 = 16'h0000;
defparam ram16s_inst_246.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_247 (
    .DO(ram16s_inst_247_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_991),
    .CLK(clk)
);

defparam ram16s_inst_247.INIT_0 = 16'h0000;
defparam ram16s_inst_247.INIT_1 = 16'h0000;
defparam ram16s_inst_247.INIT_2 = 16'h0000;
defparam ram16s_inst_247.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_248 (
    .DO(ram16s_inst_248_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_995),
    .CLK(clk)
);

defparam ram16s_inst_248.INIT_0 = 16'h0000;
defparam ram16s_inst_248.INIT_1 = 16'h0000;
defparam ram16s_inst_248.INIT_2 = 16'h0000;
defparam ram16s_inst_248.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_249 (
    .DO(ram16s_inst_249_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_999),
    .CLK(clk)
);

defparam ram16s_inst_249.INIT_0 = 16'h0000;
defparam ram16s_inst_249.INIT_1 = 16'h0000;
defparam ram16s_inst_249.INIT_2 = 16'h0000;
defparam ram16s_inst_249.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_250 (
    .DO(ram16s_inst_250_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1003),
    .CLK(clk)
);

defparam ram16s_inst_250.INIT_0 = 16'h0C00;
defparam ram16s_inst_250.INIT_1 = 16'h0000;
defparam ram16s_inst_250.INIT_2 = 16'h0000;
defparam ram16s_inst_250.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_251 (
    .DO(ram16s_inst_251_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1007),
    .CLK(clk)
);

defparam ram16s_inst_251.INIT_0 = 16'hC1C0;
defparam ram16s_inst_251.INIT_1 = 16'h0000;
defparam ram16s_inst_251.INIT_2 = 16'h0000;
defparam ram16s_inst_251.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_252 (
    .DO(ram16s_inst_252_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1011),
    .CLK(clk)
);

defparam ram16s_inst_252.INIT_0 = 16'h0384;
defparam ram16s_inst_252.INIT_1 = 16'h0000;
defparam ram16s_inst_252.INIT_2 = 16'h0000;
defparam ram16s_inst_252.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_253 (
    .DO(ram16s_inst_253_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1015),
    .CLK(clk)
);

defparam ram16s_inst_253.INIT_0 = 16'h0000;
defparam ram16s_inst_253.INIT_1 = 16'h0000;
defparam ram16s_inst_253.INIT_2 = 16'h0000;
defparam ram16s_inst_253.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_254 (
    .DO(ram16s_inst_254_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1019),
    .CLK(clk)
);

defparam ram16s_inst_254.INIT_0 = 16'h0000;
defparam ram16s_inst_254.INIT_1 = 16'h0000;
defparam ram16s_inst_254.INIT_2 = 16'h0000;
defparam ram16s_inst_254.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_255 (
    .DO(ram16s_inst_255_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1023),
    .CLK(clk)
);

defparam ram16s_inst_255.INIT_0 = 16'h0C00;
defparam ram16s_inst_255.INIT_1 = 16'h0000;
defparam ram16s_inst_255.INIT_2 = 16'h0000;
defparam ram16s_inst_255.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_256 (
    .DO(ram16s_inst_256_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1027),
    .CLK(clk)
);

defparam ram16s_inst_256.INIT_0 = 16'hC7E0;
defparam ram16s_inst_256.INIT_1 = 16'h0000;
defparam ram16s_inst_256.INIT_2 = 16'h0000;
defparam ram16s_inst_256.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_257 (
    .DO(ram16s_inst_257_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1031),
    .CLK(clk)
);

defparam ram16s_inst_257.INIT_0 = 16'h0FE7;
defparam ram16s_inst_257.INIT_1 = 16'h0000;
defparam ram16s_inst_257.INIT_2 = 16'h0000;
defparam ram16s_inst_257.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_258 (
    .DO(ram16s_inst_258_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1035),
    .CLK(clk)
);

defparam ram16s_inst_258.INIT_0 = 16'h0000;
defparam ram16s_inst_258.INIT_1 = 16'h0000;
defparam ram16s_inst_258.INIT_2 = 16'h0000;
defparam ram16s_inst_258.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_259 (
    .DO(ram16s_inst_259_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1039),
    .CLK(clk)
);

defparam ram16s_inst_259.INIT_0 = 16'h0000;
defparam ram16s_inst_259.INIT_1 = 16'h0000;
defparam ram16s_inst_259.INIT_2 = 16'h0000;
defparam ram16s_inst_259.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_260 (
    .DO(ram16s_inst_260_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1043),
    .CLK(clk)
);

defparam ram16s_inst_260.INIT_0 = 16'h0C00;
defparam ram16s_inst_260.INIT_1 = 16'h0000;
defparam ram16s_inst_260.INIT_2 = 16'h0000;
defparam ram16s_inst_260.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_261 (
    .DO(ram16s_inst_261_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1047),
    .CLK(clk)
);

defparam ram16s_inst_261.INIT_0 = 16'hCC30;
defparam ram16s_inst_261.INIT_1 = 16'h0000;
defparam ram16s_inst_261.INIT_2 = 16'h0000;
defparam ram16s_inst_261.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_262 (
    .DO(ram16s_inst_262_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1051),
    .CLK(clk)
);

defparam ram16s_inst_262.INIT_0 = 16'h0C20;
defparam ram16s_inst_262.INIT_1 = 16'h0000;
defparam ram16s_inst_262.INIT_2 = 16'h0000;
defparam ram16s_inst_262.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_263 (
    .DO(ram16s_inst_263_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1055),
    .CLK(clk)
);

defparam ram16s_inst_263.INIT_0 = 16'h0000;
defparam ram16s_inst_263.INIT_1 = 16'h0000;
defparam ram16s_inst_263.INIT_2 = 16'h0000;
defparam ram16s_inst_263.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_264 (
    .DO(ram16s_inst_264_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1059),
    .CLK(clk)
);

defparam ram16s_inst_264.INIT_0 = 16'h0000;
defparam ram16s_inst_264.INIT_1 = 16'h0000;
defparam ram16s_inst_264.INIT_2 = 16'h0000;
defparam ram16s_inst_264.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_265 (
    .DO(ram16s_inst_265_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1063),
    .CLK(clk)
);

defparam ram16s_inst_265.INIT_0 = 16'h0C00;
defparam ram16s_inst_265.INIT_1 = 16'h0000;
defparam ram16s_inst_265.INIT_2 = 16'h0000;
defparam ram16s_inst_265.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_266 (
    .DO(ram16s_inst_266_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1067),
    .CLK(clk)
);

defparam ram16s_inst_266.INIT_0 = 16'hCC10;
defparam ram16s_inst_266.INIT_1 = 16'h0000;
defparam ram16s_inst_266.INIT_2 = 16'h0000;
defparam ram16s_inst_266.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_267 (
    .DO(ram16s_inst_267_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1071),
    .CLK(clk)
);

defparam ram16s_inst_267.INIT_0 = 16'h0FF0;
defparam ram16s_inst_267.INIT_1 = 16'h0000;
defparam ram16s_inst_267.INIT_2 = 16'h0000;
defparam ram16s_inst_267.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_268 (
    .DO(ram16s_inst_268_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1075),
    .CLK(clk)
);

defparam ram16s_inst_268.INIT_0 = 16'h0000;
defparam ram16s_inst_268.INIT_1 = 16'h0000;
defparam ram16s_inst_268.INIT_2 = 16'h0000;
defparam ram16s_inst_268.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_269 (
    .DO(ram16s_inst_269_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1079),
    .CLK(clk)
);

defparam ram16s_inst_269.INIT_0 = 16'h0000;
defparam ram16s_inst_269.INIT_1 = 16'h0000;
defparam ram16s_inst_269.INIT_2 = 16'h0000;
defparam ram16s_inst_269.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_270 (
    .DO(ram16s_inst_270_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1083),
    .CLK(clk)
);

defparam ram16s_inst_270.INIT_0 = 16'h0C00;
defparam ram16s_inst_270.INIT_1 = 16'h0000;
defparam ram16s_inst_270.INIT_2 = 16'h0000;
defparam ram16s_inst_270.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_271 (
    .DO(ram16s_inst_271_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1087),
    .CLK(clk)
);

defparam ram16s_inst_271.INIT_0 = 16'hCC10;
defparam ram16s_inst_271.INIT_1 = 16'h0000;
defparam ram16s_inst_271.INIT_2 = 16'h0000;
defparam ram16s_inst_271.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_272 (
    .DO(ram16s_inst_272_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1091),
    .CLK(clk)
);

defparam ram16s_inst_272.INIT_0 = 16'h0030;
defparam ram16s_inst_272.INIT_1 = 16'h0000;
defparam ram16s_inst_272.INIT_2 = 16'h0000;
defparam ram16s_inst_272.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_273 (
    .DO(ram16s_inst_273_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1095),
    .CLK(clk)
);

defparam ram16s_inst_273.INIT_0 = 16'h0000;
defparam ram16s_inst_273.INIT_1 = 16'h0000;
defparam ram16s_inst_273.INIT_2 = 16'h0000;
defparam ram16s_inst_273.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_274 (
    .DO(ram16s_inst_274_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1099),
    .CLK(clk)
);

defparam ram16s_inst_274.INIT_0 = 16'h0000;
defparam ram16s_inst_274.INIT_1 = 16'h0000;
defparam ram16s_inst_274.INIT_2 = 16'h0000;
defparam ram16s_inst_274.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_275 (
    .DO(ram16s_inst_275_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1103),
    .CLK(clk)
);

defparam ram16s_inst_275.INIT_0 = 16'h1800;
defparam ram16s_inst_275.INIT_1 = 16'h0000;
defparam ram16s_inst_275.INIT_2 = 16'h0000;
defparam ram16s_inst_275.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_276 (
    .DO(ram16s_inst_276_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1107),
    .CLK(clk)
);

defparam ram16s_inst_276.INIT_0 = 16'hCC34;
defparam ram16s_inst_276.INIT_1 = 16'h0000;
defparam ram16s_inst_276.INIT_2 = 16'h0000;
defparam ram16s_inst_276.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_277 (
    .DO(ram16s_inst_277_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1111),
    .CLK(clk)
);

defparam ram16s_inst_277.INIT_0 = 16'h0060;
defparam ram16s_inst_277.INIT_1 = 16'h0000;
defparam ram16s_inst_277.INIT_2 = 16'h0000;
defparam ram16s_inst_277.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_278 (
    .DO(ram16s_inst_278_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1115),
    .CLK(clk)
);

defparam ram16s_inst_278.INIT_0 = 16'h0000;
defparam ram16s_inst_278.INIT_1 = 16'h0000;
defparam ram16s_inst_278.INIT_2 = 16'h0000;
defparam ram16s_inst_278.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_279 (
    .DO(ram16s_inst_279_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1119),
    .CLK(clk)
);

defparam ram16s_inst_279.INIT_0 = 16'h0000;
defparam ram16s_inst_279.INIT_1 = 16'h0000;
defparam ram16s_inst_279.INIT_2 = 16'h0000;
defparam ram16s_inst_279.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_280 (
    .DO(ram16s_inst_280_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1123),
    .CLK(clk)
);

defparam ram16s_inst_280.INIT_0 = 16'hF000;
defparam ram16s_inst_280.INIT_1 = 16'h0000;
defparam ram16s_inst_280.INIT_2 = 16'h0000;
defparam ram16s_inst_280.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_281 (
    .DO(ram16s_inst_281_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1127),
    .CLK(clk)
);

defparam ram16s_inst_281.INIT_0 = 16'hC7E7;
defparam ram16s_inst_281.INIT_1 = 16'h0000;
defparam ram16s_inst_281.INIT_2 = 16'h0000;
defparam ram16s_inst_281.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_282 (
    .DO(ram16s_inst_282_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1131),
    .CLK(clk)
);

defparam ram16s_inst_282.INIT_0 = 16'h0FE0;
defparam ram16s_inst_282.INIT_1 = 16'h0000;
defparam ram16s_inst_282.INIT_2 = 16'h0000;
defparam ram16s_inst_282.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_283 (
    .DO(ram16s_inst_283_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1135),
    .CLK(clk)
);

defparam ram16s_inst_283.INIT_0 = 16'h0000;
defparam ram16s_inst_283.INIT_1 = 16'h0000;
defparam ram16s_inst_283.INIT_2 = 16'h0000;
defparam ram16s_inst_283.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_284 (
    .DO(ram16s_inst_284_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1139),
    .CLK(clk)
);

defparam ram16s_inst_284.INIT_0 = 16'h0000;
defparam ram16s_inst_284.INIT_1 = 16'h0000;
defparam ram16s_inst_284.INIT_2 = 16'h0000;
defparam ram16s_inst_284.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_285 (
    .DO(ram16s_inst_285_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1143),
    .CLK(clk)
);

defparam ram16s_inst_285.INIT_0 = 16'hC000;
defparam ram16s_inst_285.INIT_1 = 16'h0000;
defparam ram16s_inst_285.INIT_2 = 16'h0000;
defparam ram16s_inst_285.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_286 (
    .DO(ram16s_inst_286_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1147),
    .CLK(clk)
);

defparam ram16s_inst_286.INIT_0 = 16'hC1C1;
defparam ram16s_inst_286.INIT_1 = 16'h0000;
defparam ram16s_inst_286.INIT_2 = 16'h0000;
defparam ram16s_inst_286.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_287 (
    .DO(ram16s_inst_287_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1151),
    .CLK(clk)
);

defparam ram16s_inst_287.INIT_0 = 16'h0380;
defparam ram16s_inst_287.INIT_1 = 16'h0000;
defparam ram16s_inst_287.INIT_2 = 16'h0000;
defparam ram16s_inst_287.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_288 (
    .DO(ram16s_inst_288_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1155),
    .CLK(clk)
);

defparam ram16s_inst_288.INIT_0 = 16'h0000;
defparam ram16s_inst_288.INIT_1 = 16'h0000;
defparam ram16s_inst_288.INIT_2 = 16'h0000;
defparam ram16s_inst_288.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_289 (
    .DO(ram16s_inst_289_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1159),
    .CLK(clk)
);

defparam ram16s_inst_289.INIT_0 = 16'h0000;
defparam ram16s_inst_289.INIT_1 = 16'h0000;
defparam ram16s_inst_289.INIT_2 = 16'h0000;
defparam ram16s_inst_289.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_290 (
    .DO(ram16s_inst_290_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1163),
    .CLK(clk)
);

defparam ram16s_inst_290.INIT_0 = 16'h0000;
defparam ram16s_inst_290.INIT_1 = 16'h0000;
defparam ram16s_inst_290.INIT_2 = 16'h0000;
defparam ram16s_inst_290.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_291 (
    .DO(ram16s_inst_291_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1167),
    .CLK(clk)
);

defparam ram16s_inst_291.INIT_0 = 16'h0000;
defparam ram16s_inst_291.INIT_1 = 16'h0000;
defparam ram16s_inst_291.INIT_2 = 16'h0000;
defparam ram16s_inst_291.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_292 (
    .DO(ram16s_inst_292_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1171),
    .CLK(clk)
);

defparam ram16s_inst_292.INIT_0 = 16'h0000;
defparam ram16s_inst_292.INIT_1 = 16'h0000;
defparam ram16s_inst_292.INIT_2 = 16'h0000;
defparam ram16s_inst_292.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_293 (
    .DO(ram16s_inst_293_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1175),
    .CLK(clk)
);

defparam ram16s_inst_293.INIT_0 = 16'h0000;
defparam ram16s_inst_293.INIT_1 = 16'h0000;
defparam ram16s_inst_293.INIT_2 = 16'h0000;
defparam ram16s_inst_293.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_294 (
    .DO(ram16s_inst_294_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1179),
    .CLK(clk)
);

defparam ram16s_inst_294.INIT_0 = 16'h0000;
defparam ram16s_inst_294.INIT_1 = 16'h0000;
defparam ram16s_inst_294.INIT_2 = 16'h0000;
defparam ram16s_inst_294.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_295 (
    .DO(ram16s_inst_295_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1183),
    .CLK(clk)
);

defparam ram16s_inst_295.INIT_0 = 16'h0000;
defparam ram16s_inst_295.INIT_1 = 16'h0000;
defparam ram16s_inst_295.INIT_2 = 16'h0000;
defparam ram16s_inst_295.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_296 (
    .DO(ram16s_inst_296_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1187),
    .CLK(clk)
);

defparam ram16s_inst_296.INIT_0 = 16'h0000;
defparam ram16s_inst_296.INIT_1 = 16'h0000;
defparam ram16s_inst_296.INIT_2 = 16'h0000;
defparam ram16s_inst_296.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_297 (
    .DO(ram16s_inst_297_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1191),
    .CLK(clk)
);

defparam ram16s_inst_297.INIT_0 = 16'h0000;
defparam ram16s_inst_297.INIT_1 = 16'h0000;
defparam ram16s_inst_297.INIT_2 = 16'h0000;
defparam ram16s_inst_297.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_298 (
    .DO(ram16s_inst_298_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1195),
    .CLK(clk)
);

defparam ram16s_inst_298.INIT_0 = 16'h0000;
defparam ram16s_inst_298.INIT_1 = 16'h0000;
defparam ram16s_inst_298.INIT_2 = 16'h0000;
defparam ram16s_inst_298.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_299 (
    .DO(ram16s_inst_299_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1199),
    .CLK(clk)
);

defparam ram16s_inst_299.INIT_0 = 16'h0000;
defparam ram16s_inst_299.INIT_1 = 16'h0000;
defparam ram16s_inst_299.INIT_2 = 16'h0000;
defparam ram16s_inst_299.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_300 (
    .DO(ram16s_inst_300_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1203),
    .CLK(clk)
);

defparam ram16s_inst_300.INIT_0 = 16'h0000;
defparam ram16s_inst_300.INIT_1 = 16'h0000;
defparam ram16s_inst_300.INIT_2 = 16'h0000;
defparam ram16s_inst_300.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_301 (
    .DO(ram16s_inst_301_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1207),
    .CLK(clk)
);

defparam ram16s_inst_301.INIT_0 = 16'h0000;
defparam ram16s_inst_301.INIT_1 = 16'h0000;
defparam ram16s_inst_301.INIT_2 = 16'h0000;
defparam ram16s_inst_301.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_302 (
    .DO(ram16s_inst_302_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1211),
    .CLK(clk)
);

defparam ram16s_inst_302.INIT_0 = 16'h0000;
defparam ram16s_inst_302.INIT_1 = 16'h0000;
defparam ram16s_inst_302.INIT_2 = 16'h0000;
defparam ram16s_inst_302.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_303 (
    .DO(ram16s_inst_303_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1215),
    .CLK(clk)
);

defparam ram16s_inst_303.INIT_0 = 16'h0000;
defparam ram16s_inst_303.INIT_1 = 16'h0000;
defparam ram16s_inst_303.INIT_2 = 16'h0000;
defparam ram16s_inst_303.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_304 (
    .DO(ram16s_inst_304_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1219),
    .CLK(clk)
);

defparam ram16s_inst_304.INIT_0 = 16'h0000;
defparam ram16s_inst_304.INIT_1 = 16'h0000;
defparam ram16s_inst_304.INIT_2 = 16'h0000;
defparam ram16s_inst_304.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_305 (
    .DO(ram16s_inst_305_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1223),
    .CLK(clk)
);

defparam ram16s_inst_305.INIT_0 = 16'h0000;
defparam ram16s_inst_305.INIT_1 = 16'h0000;
defparam ram16s_inst_305.INIT_2 = 16'h0000;
defparam ram16s_inst_305.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_306 (
    .DO(ram16s_inst_306_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1227),
    .CLK(clk)
);

defparam ram16s_inst_306.INIT_0 = 16'h0000;
defparam ram16s_inst_306.INIT_1 = 16'h0000;
defparam ram16s_inst_306.INIT_2 = 16'h0000;
defparam ram16s_inst_306.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_307 (
    .DO(ram16s_inst_307_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1231),
    .CLK(clk)
);

defparam ram16s_inst_307.INIT_0 = 16'h0000;
defparam ram16s_inst_307.INIT_1 = 16'h0000;
defparam ram16s_inst_307.INIT_2 = 16'h0000;
defparam ram16s_inst_307.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_308 (
    .DO(ram16s_inst_308_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1235),
    .CLK(clk)
);

defparam ram16s_inst_308.INIT_0 = 16'h0000;
defparam ram16s_inst_308.INIT_1 = 16'h0000;
defparam ram16s_inst_308.INIT_2 = 16'h0000;
defparam ram16s_inst_308.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_309 (
    .DO(ram16s_inst_309_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1239),
    .CLK(clk)
);

defparam ram16s_inst_309.INIT_0 = 16'h0000;
defparam ram16s_inst_309.INIT_1 = 16'h0000;
defparam ram16s_inst_309.INIT_2 = 16'h0000;
defparam ram16s_inst_309.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_310 (
    .DO(ram16s_inst_310_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1243),
    .CLK(clk)
);

defparam ram16s_inst_310.INIT_0 = 16'h0000;
defparam ram16s_inst_310.INIT_1 = 16'h0000;
defparam ram16s_inst_310.INIT_2 = 16'h0000;
defparam ram16s_inst_310.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_311 (
    .DO(ram16s_inst_311_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1247),
    .CLK(clk)
);

defparam ram16s_inst_311.INIT_0 = 16'h0000;
defparam ram16s_inst_311.INIT_1 = 16'h0000;
defparam ram16s_inst_311.INIT_2 = 16'h0000;
defparam ram16s_inst_311.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_312 (
    .DO(ram16s_inst_312_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1251),
    .CLK(clk)
);

defparam ram16s_inst_312.INIT_0 = 16'h0000;
defparam ram16s_inst_312.INIT_1 = 16'h0000;
defparam ram16s_inst_312.INIT_2 = 16'h0000;
defparam ram16s_inst_312.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_313 (
    .DO(ram16s_inst_313_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1255),
    .CLK(clk)
);

defparam ram16s_inst_313.INIT_0 = 16'h0000;
defparam ram16s_inst_313.INIT_1 = 16'h0000;
defparam ram16s_inst_313.INIT_2 = 16'h0000;
defparam ram16s_inst_313.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_314 (
    .DO(ram16s_inst_314_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1259),
    .CLK(clk)
);

defparam ram16s_inst_314.INIT_0 = 16'h0000;
defparam ram16s_inst_314.INIT_1 = 16'h0000;
defparam ram16s_inst_314.INIT_2 = 16'h0000;
defparam ram16s_inst_314.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_315 (
    .DO(ram16s_inst_315_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1263),
    .CLK(clk)
);

defparam ram16s_inst_315.INIT_0 = 16'h0000;
defparam ram16s_inst_315.INIT_1 = 16'h0000;
defparam ram16s_inst_315.INIT_2 = 16'h0000;
defparam ram16s_inst_315.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_316 (
    .DO(ram16s_inst_316_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1267),
    .CLK(clk)
);

defparam ram16s_inst_316.INIT_0 = 16'h0000;
defparam ram16s_inst_316.INIT_1 = 16'h0000;
defparam ram16s_inst_316.INIT_2 = 16'h0000;
defparam ram16s_inst_316.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_317 (
    .DO(ram16s_inst_317_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1271),
    .CLK(clk)
);

defparam ram16s_inst_317.INIT_0 = 16'h0000;
defparam ram16s_inst_317.INIT_1 = 16'h0000;
defparam ram16s_inst_317.INIT_2 = 16'h0000;
defparam ram16s_inst_317.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_318 (
    .DO(ram16s_inst_318_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1275),
    .CLK(clk)
);

defparam ram16s_inst_318.INIT_0 = 16'h0000;
defparam ram16s_inst_318.INIT_1 = 16'h0000;
defparam ram16s_inst_318.INIT_2 = 16'h0000;
defparam ram16s_inst_318.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_319 (
    .DO(ram16s_inst_319_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1279),
    .CLK(clk)
);

defparam ram16s_inst_319.INIT_0 = 16'h0000;
defparam ram16s_inst_319.INIT_1 = 16'h0000;
defparam ram16s_inst_319.INIT_2 = 16'h0000;
defparam ram16s_inst_319.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_320 (
    .DO(ram16s_inst_320_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1283),
    .CLK(clk)
);

defparam ram16s_inst_320.INIT_0 = 16'h0000;
defparam ram16s_inst_320.INIT_1 = 16'h0000;
defparam ram16s_inst_320.INIT_2 = 16'h0000;
defparam ram16s_inst_320.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_321 (
    .DO(ram16s_inst_321_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1287),
    .CLK(clk)
);

defparam ram16s_inst_321.INIT_0 = 16'h0000;
defparam ram16s_inst_321.INIT_1 = 16'h0000;
defparam ram16s_inst_321.INIT_2 = 16'h0000;
defparam ram16s_inst_321.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_322 (
    .DO(ram16s_inst_322_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1291),
    .CLK(clk)
);

defparam ram16s_inst_322.INIT_0 = 16'h0000;
defparam ram16s_inst_322.INIT_1 = 16'h0000;
defparam ram16s_inst_322.INIT_2 = 16'h0000;
defparam ram16s_inst_322.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_323 (
    .DO(ram16s_inst_323_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1295),
    .CLK(clk)
);

defparam ram16s_inst_323.INIT_0 = 16'h0000;
defparam ram16s_inst_323.INIT_1 = 16'h0000;
defparam ram16s_inst_323.INIT_2 = 16'h0000;
defparam ram16s_inst_323.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_324 (
    .DO(ram16s_inst_324_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1299),
    .CLK(clk)
);

defparam ram16s_inst_324.INIT_0 = 16'h0000;
defparam ram16s_inst_324.INIT_1 = 16'h0000;
defparam ram16s_inst_324.INIT_2 = 16'h0000;
defparam ram16s_inst_324.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_325 (
    .DO(ram16s_inst_325_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1303),
    .CLK(clk)
);

defparam ram16s_inst_325.INIT_0 = 16'h0000;
defparam ram16s_inst_325.INIT_1 = 16'h0000;
defparam ram16s_inst_325.INIT_2 = 16'h0000;
defparam ram16s_inst_325.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_326 (
    .DO(ram16s_inst_326_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1307),
    .CLK(clk)
);

defparam ram16s_inst_326.INIT_0 = 16'h0000;
defparam ram16s_inst_326.INIT_1 = 16'h0000;
defparam ram16s_inst_326.INIT_2 = 16'h0000;
defparam ram16s_inst_326.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_327 (
    .DO(ram16s_inst_327_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1311),
    .CLK(clk)
);

defparam ram16s_inst_327.INIT_0 = 16'h0000;
defparam ram16s_inst_327.INIT_1 = 16'h0000;
defparam ram16s_inst_327.INIT_2 = 16'h0000;
defparam ram16s_inst_327.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_328 (
    .DO(ram16s_inst_328_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1315),
    .CLK(clk)
);

defparam ram16s_inst_328.INIT_0 = 16'h0000;
defparam ram16s_inst_328.INIT_1 = 16'h0000;
defparam ram16s_inst_328.INIT_2 = 16'h0000;
defparam ram16s_inst_328.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_329 (
    .DO(ram16s_inst_329_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1319),
    .CLK(clk)
);

defparam ram16s_inst_329.INIT_0 = 16'h0000;
defparam ram16s_inst_329.INIT_1 = 16'h0000;
defparam ram16s_inst_329.INIT_2 = 16'h0000;
defparam ram16s_inst_329.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_330 (
    .DO(ram16s_inst_330_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1323),
    .CLK(clk)
);

defparam ram16s_inst_330.INIT_0 = 16'h0000;
defparam ram16s_inst_330.INIT_1 = 16'h0000;
defparam ram16s_inst_330.INIT_2 = 16'h0000;
defparam ram16s_inst_330.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_331 (
    .DO(ram16s_inst_331_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1327),
    .CLK(clk)
);

defparam ram16s_inst_331.INIT_0 = 16'h0000;
defparam ram16s_inst_331.INIT_1 = 16'h0000;
defparam ram16s_inst_331.INIT_2 = 16'h0000;
defparam ram16s_inst_331.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_332 (
    .DO(ram16s_inst_332_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1331),
    .CLK(clk)
);

defparam ram16s_inst_332.INIT_0 = 16'h0000;
defparam ram16s_inst_332.INIT_1 = 16'h0000;
defparam ram16s_inst_332.INIT_2 = 16'h0000;
defparam ram16s_inst_332.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_333 (
    .DO(ram16s_inst_333_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1335),
    .CLK(clk)
);

defparam ram16s_inst_333.INIT_0 = 16'h0000;
defparam ram16s_inst_333.INIT_1 = 16'h0000;
defparam ram16s_inst_333.INIT_2 = 16'h0000;
defparam ram16s_inst_333.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_334 (
    .DO(ram16s_inst_334_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1339),
    .CLK(clk)
);

defparam ram16s_inst_334.INIT_0 = 16'h0000;
defparam ram16s_inst_334.INIT_1 = 16'h0000;
defparam ram16s_inst_334.INIT_2 = 16'h0000;
defparam ram16s_inst_334.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_335 (
    .DO(ram16s_inst_335_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1343),
    .CLK(clk)
);

defparam ram16s_inst_335.INIT_0 = 16'h0000;
defparam ram16s_inst_335.INIT_1 = 16'h0000;
defparam ram16s_inst_335.INIT_2 = 16'h0000;
defparam ram16s_inst_335.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_336 (
    .DO(ram16s_inst_336_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1347),
    .CLK(clk)
);

defparam ram16s_inst_336.INIT_0 = 16'h0000;
defparam ram16s_inst_336.INIT_1 = 16'h0000;
defparam ram16s_inst_336.INIT_2 = 16'h0000;
defparam ram16s_inst_336.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_337 (
    .DO(ram16s_inst_337_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1351),
    .CLK(clk)
);

defparam ram16s_inst_337.INIT_0 = 16'h0000;
defparam ram16s_inst_337.INIT_1 = 16'h0000;
defparam ram16s_inst_337.INIT_2 = 16'h0000;
defparam ram16s_inst_337.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_338 (
    .DO(ram16s_inst_338_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1355),
    .CLK(clk)
);

defparam ram16s_inst_338.INIT_0 = 16'h0000;
defparam ram16s_inst_338.INIT_1 = 16'h0000;
defparam ram16s_inst_338.INIT_2 = 16'h0000;
defparam ram16s_inst_338.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_339 (
    .DO(ram16s_inst_339_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1359),
    .CLK(clk)
);

defparam ram16s_inst_339.INIT_0 = 16'h0000;
defparam ram16s_inst_339.INIT_1 = 16'h0000;
defparam ram16s_inst_339.INIT_2 = 16'h0000;
defparam ram16s_inst_339.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_340 (
    .DO(ram16s_inst_340_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1363),
    .CLK(clk)
);

defparam ram16s_inst_340.INIT_0 = 16'h0000;
defparam ram16s_inst_340.INIT_1 = 16'h0000;
defparam ram16s_inst_340.INIT_2 = 16'h0000;
defparam ram16s_inst_340.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_341 (
    .DO(ram16s_inst_341_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1367),
    .CLK(clk)
);

defparam ram16s_inst_341.INIT_0 = 16'h0000;
defparam ram16s_inst_341.INIT_1 = 16'h0000;
defparam ram16s_inst_341.INIT_2 = 16'h0000;
defparam ram16s_inst_341.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_342 (
    .DO(ram16s_inst_342_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1371),
    .CLK(clk)
);

defparam ram16s_inst_342.INIT_0 = 16'h0000;
defparam ram16s_inst_342.INIT_1 = 16'h0000;
defparam ram16s_inst_342.INIT_2 = 16'h0000;
defparam ram16s_inst_342.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_343 (
    .DO(ram16s_inst_343_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1375),
    .CLK(clk)
);

defparam ram16s_inst_343.INIT_0 = 16'h0000;
defparam ram16s_inst_343.INIT_1 = 16'h0000;
defparam ram16s_inst_343.INIT_2 = 16'h0000;
defparam ram16s_inst_343.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_344 (
    .DO(ram16s_inst_344_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1379),
    .CLK(clk)
);

defparam ram16s_inst_344.INIT_0 = 16'h0000;
defparam ram16s_inst_344.INIT_1 = 16'h0000;
defparam ram16s_inst_344.INIT_2 = 16'h0000;
defparam ram16s_inst_344.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_345 (
    .DO(ram16s_inst_345_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1383),
    .CLK(clk)
);

defparam ram16s_inst_345.INIT_0 = 16'h0000;
defparam ram16s_inst_345.INIT_1 = 16'h0000;
defparam ram16s_inst_345.INIT_2 = 16'hFE00;
defparam ram16s_inst_345.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_346 (
    .DO(ram16s_inst_346_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1387),
    .CLK(clk)
);

defparam ram16s_inst_346.INIT_0 = 16'h0000;
defparam ram16s_inst_346.INIT_1 = 16'h0000;
defparam ram16s_inst_346.INIT_2 = 16'h87F0;
defparam ram16s_inst_346.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_347 (
    .DO(ram16s_inst_347_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1391),
    .CLK(clk)
);

defparam ram16s_inst_347.INIT_0 = 16'h0000;
defparam ram16s_inst_347.INIT_1 = 16'h0000;
defparam ram16s_inst_347.INIT_2 = 16'hFC3F;
defparam ram16s_inst_347.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_348 (
    .DO(ram16s_inst_348_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1395),
    .CLK(clk)
);

defparam ram16s_inst_348.INIT_0 = 16'h0000;
defparam ram16s_inst_348.INIT_1 = 16'h0000;
defparam ram16s_inst_348.INIT_2 = 16'h07F1;
defparam ram16s_inst_348.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_349 (
    .DO(ram16s_inst_349_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1399),
    .CLK(clk)
);

defparam ram16s_inst_349.INIT_0 = 16'h0000;
defparam ram16s_inst_349.INIT_1 = 16'h0000;
defparam ram16s_inst_349.INIT_2 = 16'h0000;
defparam ram16s_inst_349.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_350 (
    .DO(ram16s_inst_350_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1403),
    .CLK(clk)
);

defparam ram16s_inst_350.INIT_0 = 16'h0000;
defparam ram16s_inst_350.INIT_1 = 16'h0000;
defparam ram16s_inst_350.INIT_2 = 16'hFE00;
defparam ram16s_inst_350.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_351 (
    .DO(ram16s_inst_351_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1407),
    .CLK(clk)
);

defparam ram16s_inst_351.INIT_0 = 16'h0000;
defparam ram16s_inst_351.INIT_1 = 16'h0000;
defparam ram16s_inst_351.INIT_2 = 16'h87F0;
defparam ram16s_inst_351.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_352 (
    .DO(ram16s_inst_352_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1411),
    .CLK(clk)
);

defparam ram16s_inst_352.INIT_0 = 16'h0000;
defparam ram16s_inst_352.INIT_1 = 16'h0000;
defparam ram16s_inst_352.INIT_2 = 16'hFC3F;
defparam ram16s_inst_352.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_353 (
    .DO(ram16s_inst_353_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1415),
    .CLK(clk)
);

defparam ram16s_inst_353.INIT_0 = 16'h0000;
defparam ram16s_inst_353.INIT_1 = 16'h0000;
defparam ram16s_inst_353.INIT_2 = 16'h07F1;
defparam ram16s_inst_353.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_354 (
    .DO(ram16s_inst_354_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1419),
    .CLK(clk)
);

defparam ram16s_inst_354.INIT_0 = 16'h0000;
defparam ram16s_inst_354.INIT_1 = 16'h0000;
defparam ram16s_inst_354.INIT_2 = 16'h0000;
defparam ram16s_inst_354.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_355 (
    .DO(ram16s_inst_355_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1423),
    .CLK(clk)
);

defparam ram16s_inst_355.INIT_0 = 16'h0000;
defparam ram16s_inst_355.INIT_1 = 16'h0000;
defparam ram16s_inst_355.INIT_2 = 16'hFE00;
defparam ram16s_inst_355.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_356 (
    .DO(ram16s_inst_356_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1427),
    .CLK(clk)
);

defparam ram16s_inst_356.INIT_0 = 16'h0000;
defparam ram16s_inst_356.INIT_1 = 16'h0000;
defparam ram16s_inst_356.INIT_2 = 16'h87F0;
defparam ram16s_inst_356.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_357 (
    .DO(ram16s_inst_357_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1431),
    .CLK(clk)
);

defparam ram16s_inst_357.INIT_0 = 16'h0000;
defparam ram16s_inst_357.INIT_1 = 16'h0000;
defparam ram16s_inst_357.INIT_2 = 16'hFC3F;
defparam ram16s_inst_357.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_358 (
    .DO(ram16s_inst_358_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1435),
    .CLK(clk)
);

defparam ram16s_inst_358.INIT_0 = 16'h0000;
defparam ram16s_inst_358.INIT_1 = 16'h0000;
defparam ram16s_inst_358.INIT_2 = 16'h07F1;
defparam ram16s_inst_358.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_359 (
    .DO(ram16s_inst_359_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1439),
    .CLK(clk)
);

defparam ram16s_inst_359.INIT_0 = 16'h0000;
defparam ram16s_inst_359.INIT_1 = 16'h0000;
defparam ram16s_inst_359.INIT_2 = 16'h0000;
defparam ram16s_inst_359.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_360 (
    .DO(ram16s_inst_360_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1443),
    .CLK(clk)
);

defparam ram16s_inst_360.INIT_0 = 16'h0000;
defparam ram16s_inst_360.INIT_1 = 16'h0000;
defparam ram16s_inst_360.INIT_2 = 16'hFE00;
defparam ram16s_inst_360.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_361 (
    .DO(ram16s_inst_361_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1447),
    .CLK(clk)
);

defparam ram16s_inst_361.INIT_0 = 16'h0000;
defparam ram16s_inst_361.INIT_1 = 16'h0000;
defparam ram16s_inst_361.INIT_2 = 16'h87F0;
defparam ram16s_inst_361.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_362 (
    .DO(ram16s_inst_362_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1451),
    .CLK(clk)
);

defparam ram16s_inst_362.INIT_0 = 16'h0000;
defparam ram16s_inst_362.INIT_1 = 16'h0000;
defparam ram16s_inst_362.INIT_2 = 16'hFC3F;
defparam ram16s_inst_362.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_363 (
    .DO(ram16s_inst_363_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1455),
    .CLK(clk)
);

defparam ram16s_inst_363.INIT_0 = 16'h0000;
defparam ram16s_inst_363.INIT_1 = 16'h0000;
defparam ram16s_inst_363.INIT_2 = 16'h07F1;
defparam ram16s_inst_363.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_364 (
    .DO(ram16s_inst_364_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1459),
    .CLK(clk)
);

defparam ram16s_inst_364.INIT_0 = 16'h0000;
defparam ram16s_inst_364.INIT_1 = 16'h0000;
defparam ram16s_inst_364.INIT_2 = 16'h0000;
defparam ram16s_inst_364.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_365 (
    .DO(ram16s_inst_365_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1463),
    .CLK(clk)
);

defparam ram16s_inst_365.INIT_0 = 16'h0000;
defparam ram16s_inst_365.INIT_1 = 16'h0000;
defparam ram16s_inst_365.INIT_2 = 16'hFE00;
defparam ram16s_inst_365.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_366 (
    .DO(ram16s_inst_366_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1467),
    .CLK(clk)
);

defparam ram16s_inst_366.INIT_0 = 16'h0000;
defparam ram16s_inst_366.INIT_1 = 16'h0000;
defparam ram16s_inst_366.INIT_2 = 16'h87F0;
defparam ram16s_inst_366.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_367 (
    .DO(ram16s_inst_367_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1471),
    .CLK(clk)
);

defparam ram16s_inst_367.INIT_0 = 16'h0000;
defparam ram16s_inst_367.INIT_1 = 16'h0000;
defparam ram16s_inst_367.INIT_2 = 16'hFC3F;
defparam ram16s_inst_367.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_368 (
    .DO(ram16s_inst_368_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1475),
    .CLK(clk)
);

defparam ram16s_inst_368.INIT_0 = 16'h0000;
defparam ram16s_inst_368.INIT_1 = 16'h0000;
defparam ram16s_inst_368.INIT_2 = 16'h07F1;
defparam ram16s_inst_368.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_369 (
    .DO(ram16s_inst_369_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1479),
    .CLK(clk)
);

defparam ram16s_inst_369.INIT_0 = 16'h0000;
defparam ram16s_inst_369.INIT_1 = 16'h0000;
defparam ram16s_inst_369.INIT_2 = 16'h0000;
defparam ram16s_inst_369.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_370 (
    .DO(ram16s_inst_370_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1483),
    .CLK(clk)
);

defparam ram16s_inst_370.INIT_0 = 16'h0000;
defparam ram16s_inst_370.INIT_1 = 16'h0000;
defparam ram16s_inst_370.INIT_2 = 16'hFE00;
defparam ram16s_inst_370.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_371 (
    .DO(ram16s_inst_371_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1487),
    .CLK(clk)
);

defparam ram16s_inst_371.INIT_0 = 16'h0000;
defparam ram16s_inst_371.INIT_1 = 16'h0000;
defparam ram16s_inst_371.INIT_2 = 16'h87F0;
defparam ram16s_inst_371.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_372 (
    .DO(ram16s_inst_372_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1491),
    .CLK(clk)
);

defparam ram16s_inst_372.INIT_0 = 16'h0000;
defparam ram16s_inst_372.INIT_1 = 16'h0000;
defparam ram16s_inst_372.INIT_2 = 16'hFC3F;
defparam ram16s_inst_372.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_373 (
    .DO(ram16s_inst_373_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1495),
    .CLK(clk)
);

defparam ram16s_inst_373.INIT_0 = 16'h0000;
defparam ram16s_inst_373.INIT_1 = 16'h0000;
defparam ram16s_inst_373.INIT_2 = 16'h07F1;
defparam ram16s_inst_373.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_374 (
    .DO(ram16s_inst_374_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1499),
    .CLK(clk)
);

defparam ram16s_inst_374.INIT_0 = 16'h0000;
defparam ram16s_inst_374.INIT_1 = 16'h0000;
defparam ram16s_inst_374.INIT_2 = 16'h0000;
defparam ram16s_inst_374.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_375 (
    .DO(ram16s_inst_375_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1503),
    .CLK(clk)
);

defparam ram16s_inst_375.INIT_0 = 16'h0000;
defparam ram16s_inst_375.INIT_1 = 16'h0000;
defparam ram16s_inst_375.INIT_2 = 16'hFE00;
defparam ram16s_inst_375.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_376 (
    .DO(ram16s_inst_376_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1507),
    .CLK(clk)
);

defparam ram16s_inst_376.INIT_0 = 16'h0000;
defparam ram16s_inst_376.INIT_1 = 16'h0000;
defparam ram16s_inst_376.INIT_2 = 16'h87F0;
defparam ram16s_inst_376.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_377 (
    .DO(ram16s_inst_377_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1511),
    .CLK(clk)
);

defparam ram16s_inst_377.INIT_0 = 16'h0000;
defparam ram16s_inst_377.INIT_1 = 16'h0000;
defparam ram16s_inst_377.INIT_2 = 16'hFC3F;
defparam ram16s_inst_377.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_378 (
    .DO(ram16s_inst_378_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1515),
    .CLK(clk)
);

defparam ram16s_inst_378.INIT_0 = 16'h0000;
defparam ram16s_inst_378.INIT_1 = 16'h0000;
defparam ram16s_inst_378.INIT_2 = 16'h07F1;
defparam ram16s_inst_378.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_379 (
    .DO(ram16s_inst_379_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1519),
    .CLK(clk)
);

defparam ram16s_inst_379.INIT_0 = 16'h0000;
defparam ram16s_inst_379.INIT_1 = 16'h0000;
defparam ram16s_inst_379.INIT_2 = 16'h0000;
defparam ram16s_inst_379.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_380 (
    .DO(ram16s_inst_380_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1523),
    .CLK(clk)
);

defparam ram16s_inst_380.INIT_0 = 16'h0000;
defparam ram16s_inst_380.INIT_1 = 16'h0000;
defparam ram16s_inst_380.INIT_2 = 16'hFE00;
defparam ram16s_inst_380.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_381 (
    .DO(ram16s_inst_381_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1527),
    .CLK(clk)
);

defparam ram16s_inst_381.INIT_0 = 16'h0000;
defparam ram16s_inst_381.INIT_1 = 16'h0000;
defparam ram16s_inst_381.INIT_2 = 16'h87F0;
defparam ram16s_inst_381.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_382 (
    .DO(ram16s_inst_382_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1531),
    .CLK(clk)
);

defparam ram16s_inst_382.INIT_0 = 16'h0000;
defparam ram16s_inst_382.INIT_1 = 16'h0000;
defparam ram16s_inst_382.INIT_2 = 16'hFC3F;
defparam ram16s_inst_382.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_383 (
    .DO(ram16s_inst_383_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1535),
    .CLK(clk)
);

defparam ram16s_inst_383.INIT_0 = 16'h0000;
defparam ram16s_inst_383.INIT_1 = 16'h0000;
defparam ram16s_inst_383.INIT_2 = 16'h07F1;
defparam ram16s_inst_383.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_384 (
    .DO(ram16s_inst_384_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1539),
    .CLK(clk)
);

defparam ram16s_inst_384.INIT_0 = 16'h0000;
defparam ram16s_inst_384.INIT_1 = 16'h0000;
defparam ram16s_inst_384.INIT_2 = 16'h0000;
defparam ram16s_inst_384.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_385 (
    .DO(ram16s_inst_385_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1543),
    .CLK(clk)
);

defparam ram16s_inst_385.INIT_0 = 16'h0000;
defparam ram16s_inst_385.INIT_1 = 16'h0000;
defparam ram16s_inst_385.INIT_2 = 16'hFE00;
defparam ram16s_inst_385.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_386 (
    .DO(ram16s_inst_386_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1547),
    .CLK(clk)
);

defparam ram16s_inst_386.INIT_0 = 16'h0000;
defparam ram16s_inst_386.INIT_1 = 16'h0000;
defparam ram16s_inst_386.INIT_2 = 16'h87F0;
defparam ram16s_inst_386.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_387 (
    .DO(ram16s_inst_387_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1551),
    .CLK(clk)
);

defparam ram16s_inst_387.INIT_0 = 16'h0000;
defparam ram16s_inst_387.INIT_1 = 16'h0000;
defparam ram16s_inst_387.INIT_2 = 16'hFC3F;
defparam ram16s_inst_387.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_388 (
    .DO(ram16s_inst_388_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1555),
    .CLK(clk)
);

defparam ram16s_inst_388.INIT_0 = 16'h0000;
defparam ram16s_inst_388.INIT_1 = 16'h0000;
defparam ram16s_inst_388.INIT_2 = 16'h07F1;
defparam ram16s_inst_388.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_389 (
    .DO(ram16s_inst_389_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1559),
    .CLK(clk)
);

defparam ram16s_inst_389.INIT_0 = 16'h0000;
defparam ram16s_inst_389.INIT_1 = 16'h0000;
defparam ram16s_inst_389.INIT_2 = 16'h0000;
defparam ram16s_inst_389.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_390 (
    .DO(ram16s_inst_390_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1563),
    .CLK(clk)
);

defparam ram16s_inst_390.INIT_0 = 16'h0000;
defparam ram16s_inst_390.INIT_1 = 16'h0000;
defparam ram16s_inst_390.INIT_2 = 16'hFE00;
defparam ram16s_inst_390.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_391 (
    .DO(ram16s_inst_391_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1567),
    .CLK(clk)
);

defparam ram16s_inst_391.INIT_0 = 16'h0000;
defparam ram16s_inst_391.INIT_1 = 16'h0000;
defparam ram16s_inst_391.INIT_2 = 16'h87F0;
defparam ram16s_inst_391.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_392 (
    .DO(ram16s_inst_392_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1571),
    .CLK(clk)
);

defparam ram16s_inst_392.INIT_0 = 16'h0000;
defparam ram16s_inst_392.INIT_1 = 16'h0000;
defparam ram16s_inst_392.INIT_2 = 16'hFC3F;
defparam ram16s_inst_392.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_393 (
    .DO(ram16s_inst_393_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1575),
    .CLK(clk)
);

defparam ram16s_inst_393.INIT_0 = 16'h0000;
defparam ram16s_inst_393.INIT_1 = 16'h0000;
defparam ram16s_inst_393.INIT_2 = 16'h07F1;
defparam ram16s_inst_393.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_394 (
    .DO(ram16s_inst_394_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1579),
    .CLK(clk)
);

defparam ram16s_inst_394.INIT_0 = 16'h0000;
defparam ram16s_inst_394.INIT_1 = 16'h0000;
defparam ram16s_inst_394.INIT_2 = 16'h0000;
defparam ram16s_inst_394.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_395 (
    .DO(ram16s_inst_395_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1583),
    .CLK(clk)
);

defparam ram16s_inst_395.INIT_0 = 16'h0000;
defparam ram16s_inst_395.INIT_1 = 16'h0000;
defparam ram16s_inst_395.INIT_2 = 16'hFE00;
defparam ram16s_inst_395.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_396 (
    .DO(ram16s_inst_396_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1587),
    .CLK(clk)
);

defparam ram16s_inst_396.INIT_0 = 16'h0000;
defparam ram16s_inst_396.INIT_1 = 16'h0000;
defparam ram16s_inst_396.INIT_2 = 16'h87F0;
defparam ram16s_inst_396.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_397 (
    .DO(ram16s_inst_397_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1591),
    .CLK(clk)
);

defparam ram16s_inst_397.INIT_0 = 16'h0000;
defparam ram16s_inst_397.INIT_1 = 16'h0000;
defparam ram16s_inst_397.INIT_2 = 16'hFC3F;
defparam ram16s_inst_397.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_398 (
    .DO(ram16s_inst_398_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1595),
    .CLK(clk)
);

defparam ram16s_inst_398.INIT_0 = 16'h0000;
defparam ram16s_inst_398.INIT_1 = 16'h0000;
defparam ram16s_inst_398.INIT_2 = 16'h07F1;
defparam ram16s_inst_398.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_399 (
    .DO(ram16s_inst_399_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1599),
    .CLK(clk)
);

defparam ram16s_inst_399.INIT_0 = 16'h0000;
defparam ram16s_inst_399.INIT_1 = 16'h0000;
defparam ram16s_inst_399.INIT_2 = 16'h0000;
defparam ram16s_inst_399.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_400 (
    .DO(ram16s_inst_400_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1603),
    .CLK(clk)
);

defparam ram16s_inst_400.INIT_0 = 16'h0000;
defparam ram16s_inst_400.INIT_1 = 16'h0000;
defparam ram16s_inst_400.INIT_2 = 16'hFE00;
defparam ram16s_inst_400.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_401 (
    .DO(ram16s_inst_401_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1607),
    .CLK(clk)
);

defparam ram16s_inst_401.INIT_0 = 16'h0000;
defparam ram16s_inst_401.INIT_1 = 16'h0000;
defparam ram16s_inst_401.INIT_2 = 16'h87F0;
defparam ram16s_inst_401.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_402 (
    .DO(ram16s_inst_402_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1611),
    .CLK(clk)
);

defparam ram16s_inst_402.INIT_0 = 16'h0000;
defparam ram16s_inst_402.INIT_1 = 16'h0000;
defparam ram16s_inst_402.INIT_2 = 16'hFC3F;
defparam ram16s_inst_402.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_403 (
    .DO(ram16s_inst_403_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1615),
    .CLK(clk)
);

defparam ram16s_inst_403.INIT_0 = 16'h0000;
defparam ram16s_inst_403.INIT_1 = 16'h0000;
defparam ram16s_inst_403.INIT_2 = 16'h07F1;
defparam ram16s_inst_403.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_404 (
    .DO(ram16s_inst_404_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1619),
    .CLK(clk)
);

defparam ram16s_inst_404.INIT_0 = 16'h0000;
defparam ram16s_inst_404.INIT_1 = 16'h0000;
defparam ram16s_inst_404.INIT_2 = 16'h0000;
defparam ram16s_inst_404.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_405 (
    .DO(ram16s_inst_405_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1623),
    .CLK(clk)
);

defparam ram16s_inst_405.INIT_0 = 16'h0000;
defparam ram16s_inst_405.INIT_1 = 16'h0000;
defparam ram16s_inst_405.INIT_2 = 16'hFE00;
defparam ram16s_inst_405.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_406 (
    .DO(ram16s_inst_406_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1627),
    .CLK(clk)
);

defparam ram16s_inst_406.INIT_0 = 16'h0000;
defparam ram16s_inst_406.INIT_1 = 16'h0000;
defparam ram16s_inst_406.INIT_2 = 16'h87F0;
defparam ram16s_inst_406.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_407 (
    .DO(ram16s_inst_407_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1631),
    .CLK(clk)
);

defparam ram16s_inst_407.INIT_0 = 16'h0000;
defparam ram16s_inst_407.INIT_1 = 16'h0000;
defparam ram16s_inst_407.INIT_2 = 16'hFC3F;
defparam ram16s_inst_407.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_408 (
    .DO(ram16s_inst_408_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1635),
    .CLK(clk)
);

defparam ram16s_inst_408.INIT_0 = 16'h0000;
defparam ram16s_inst_408.INIT_1 = 16'h0000;
defparam ram16s_inst_408.INIT_2 = 16'h07F1;
defparam ram16s_inst_408.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_409 (
    .DO(ram16s_inst_409_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1639),
    .CLK(clk)
);

defparam ram16s_inst_409.INIT_0 = 16'h0000;
defparam ram16s_inst_409.INIT_1 = 16'h0000;
defparam ram16s_inst_409.INIT_2 = 16'h0000;
defparam ram16s_inst_409.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_410 (
    .DO(ram16s_inst_410_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1643),
    .CLK(clk)
);

defparam ram16s_inst_410.INIT_0 = 16'h0000;
defparam ram16s_inst_410.INIT_1 = 16'h0000;
defparam ram16s_inst_410.INIT_2 = 16'hFE00;
defparam ram16s_inst_410.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_411 (
    .DO(ram16s_inst_411_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1647),
    .CLK(clk)
);

defparam ram16s_inst_411.INIT_0 = 16'h0000;
defparam ram16s_inst_411.INIT_1 = 16'h0000;
defparam ram16s_inst_411.INIT_2 = 16'h87F0;
defparam ram16s_inst_411.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_412 (
    .DO(ram16s_inst_412_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1651),
    .CLK(clk)
);

defparam ram16s_inst_412.INIT_0 = 16'h0000;
defparam ram16s_inst_412.INIT_1 = 16'h0000;
defparam ram16s_inst_412.INIT_2 = 16'hFC3F;
defparam ram16s_inst_412.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_413 (
    .DO(ram16s_inst_413_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1655),
    .CLK(clk)
);

defparam ram16s_inst_413.INIT_0 = 16'h0000;
defparam ram16s_inst_413.INIT_1 = 16'h0000;
defparam ram16s_inst_413.INIT_2 = 16'h07F1;
defparam ram16s_inst_413.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_414 (
    .DO(ram16s_inst_414_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1659),
    .CLK(clk)
);

defparam ram16s_inst_414.INIT_0 = 16'h0000;
defparam ram16s_inst_414.INIT_1 = 16'h0000;
defparam ram16s_inst_414.INIT_2 = 16'h0000;
defparam ram16s_inst_414.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_415 (
    .DO(ram16s_inst_415_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1663),
    .CLK(clk)
);

defparam ram16s_inst_415.INIT_0 = 16'h0000;
defparam ram16s_inst_415.INIT_1 = 16'h0000;
defparam ram16s_inst_415.INIT_2 = 16'h0000;
defparam ram16s_inst_415.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_416 (
    .DO(ram16s_inst_416_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1667),
    .CLK(clk)
);

defparam ram16s_inst_416.INIT_0 = 16'h0000;
defparam ram16s_inst_416.INIT_1 = 16'h0000;
defparam ram16s_inst_416.INIT_2 = 16'h0000;
defparam ram16s_inst_416.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_417 (
    .DO(ram16s_inst_417_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1671),
    .CLK(clk)
);

defparam ram16s_inst_417.INIT_0 = 16'h0000;
defparam ram16s_inst_417.INIT_1 = 16'h0000;
defparam ram16s_inst_417.INIT_2 = 16'h0000;
defparam ram16s_inst_417.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_418 (
    .DO(ram16s_inst_418_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1675),
    .CLK(clk)
);

defparam ram16s_inst_418.INIT_0 = 16'h0000;
defparam ram16s_inst_418.INIT_1 = 16'h0000;
defparam ram16s_inst_418.INIT_2 = 16'h0000;
defparam ram16s_inst_418.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_419 (
    .DO(ram16s_inst_419_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1679),
    .CLK(clk)
);

defparam ram16s_inst_419.INIT_0 = 16'h0000;
defparam ram16s_inst_419.INIT_1 = 16'h0000;
defparam ram16s_inst_419.INIT_2 = 16'h0000;
defparam ram16s_inst_419.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_420 (
    .DO(ram16s_inst_420_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1683),
    .CLK(clk)
);

defparam ram16s_inst_420.INIT_0 = 16'h0000;
defparam ram16s_inst_420.INIT_1 = 16'h0000;
defparam ram16s_inst_420.INIT_2 = 16'h0000;
defparam ram16s_inst_420.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_421 (
    .DO(ram16s_inst_421_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1687),
    .CLK(clk)
);

defparam ram16s_inst_421.INIT_0 = 16'h0000;
defparam ram16s_inst_421.INIT_1 = 16'h0000;
defparam ram16s_inst_421.INIT_2 = 16'h0000;
defparam ram16s_inst_421.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_422 (
    .DO(ram16s_inst_422_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1691),
    .CLK(clk)
);

defparam ram16s_inst_422.INIT_0 = 16'h0000;
defparam ram16s_inst_422.INIT_1 = 16'h0000;
defparam ram16s_inst_422.INIT_2 = 16'h0000;
defparam ram16s_inst_422.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_423 (
    .DO(ram16s_inst_423_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1695),
    .CLK(clk)
);

defparam ram16s_inst_423.INIT_0 = 16'h0000;
defparam ram16s_inst_423.INIT_1 = 16'h0000;
defparam ram16s_inst_423.INIT_2 = 16'h0000;
defparam ram16s_inst_423.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_424 (
    .DO(ram16s_inst_424_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1699),
    .CLK(clk)
);

defparam ram16s_inst_424.INIT_0 = 16'h0000;
defparam ram16s_inst_424.INIT_1 = 16'h0000;
defparam ram16s_inst_424.INIT_2 = 16'h0000;
defparam ram16s_inst_424.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_425 (
    .DO(ram16s_inst_425_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1703),
    .CLK(clk)
);

defparam ram16s_inst_425.INIT_0 = 16'h0000;
defparam ram16s_inst_425.INIT_1 = 16'h0000;
defparam ram16s_inst_425.INIT_2 = 16'h0000;
defparam ram16s_inst_425.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_426 (
    .DO(ram16s_inst_426_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1707),
    .CLK(clk)
);

defparam ram16s_inst_426.INIT_0 = 16'h0000;
defparam ram16s_inst_426.INIT_1 = 16'h0000;
defparam ram16s_inst_426.INIT_2 = 16'h0000;
defparam ram16s_inst_426.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_427 (
    .DO(ram16s_inst_427_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1711),
    .CLK(clk)
);

defparam ram16s_inst_427.INIT_0 = 16'h0000;
defparam ram16s_inst_427.INIT_1 = 16'h0000;
defparam ram16s_inst_427.INIT_2 = 16'h0000;
defparam ram16s_inst_427.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_428 (
    .DO(ram16s_inst_428_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1715),
    .CLK(clk)
);

defparam ram16s_inst_428.INIT_0 = 16'h0000;
defparam ram16s_inst_428.INIT_1 = 16'h0000;
defparam ram16s_inst_428.INIT_2 = 16'h0000;
defparam ram16s_inst_428.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_429 (
    .DO(ram16s_inst_429_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1719),
    .CLK(clk)
);

defparam ram16s_inst_429.INIT_0 = 16'h0000;
defparam ram16s_inst_429.INIT_1 = 16'h0000;
defparam ram16s_inst_429.INIT_2 = 16'h0000;
defparam ram16s_inst_429.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_430 (
    .DO(ram16s_inst_430_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1723),
    .CLK(clk)
);

defparam ram16s_inst_430.INIT_0 = 16'h0000;
defparam ram16s_inst_430.INIT_1 = 16'h0000;
defparam ram16s_inst_430.INIT_2 = 16'h0000;
defparam ram16s_inst_430.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_431 (
    .DO(ram16s_inst_431_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1727),
    .CLK(clk)
);

defparam ram16s_inst_431.INIT_0 = 16'h0000;
defparam ram16s_inst_431.INIT_1 = 16'h0000;
defparam ram16s_inst_431.INIT_2 = 16'h0000;
defparam ram16s_inst_431.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_432 (
    .DO(ram16s_inst_432_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1731),
    .CLK(clk)
);

defparam ram16s_inst_432.INIT_0 = 16'h0000;
defparam ram16s_inst_432.INIT_1 = 16'h0000;
defparam ram16s_inst_432.INIT_2 = 16'h0000;
defparam ram16s_inst_432.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_433 (
    .DO(ram16s_inst_433_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1735),
    .CLK(clk)
);

defparam ram16s_inst_433.INIT_0 = 16'h0000;
defparam ram16s_inst_433.INIT_1 = 16'h0000;
defparam ram16s_inst_433.INIT_2 = 16'h0000;
defparam ram16s_inst_433.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_434 (
    .DO(ram16s_inst_434_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1739),
    .CLK(clk)
);

defparam ram16s_inst_434.INIT_0 = 16'h0000;
defparam ram16s_inst_434.INIT_1 = 16'h0000;
defparam ram16s_inst_434.INIT_2 = 16'h0000;
defparam ram16s_inst_434.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_435 (
    .DO(ram16s_inst_435_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1743),
    .CLK(clk)
);

defparam ram16s_inst_435.INIT_0 = 16'h0000;
defparam ram16s_inst_435.INIT_1 = 16'h0000;
defparam ram16s_inst_435.INIT_2 = 16'h0000;
defparam ram16s_inst_435.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_436 (
    .DO(ram16s_inst_436_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1747),
    .CLK(clk)
);

defparam ram16s_inst_436.INIT_0 = 16'h0000;
defparam ram16s_inst_436.INIT_1 = 16'h0000;
defparam ram16s_inst_436.INIT_2 = 16'h0000;
defparam ram16s_inst_436.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_437 (
    .DO(ram16s_inst_437_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1751),
    .CLK(clk)
);

defparam ram16s_inst_437.INIT_0 = 16'h0000;
defparam ram16s_inst_437.INIT_1 = 16'h0000;
defparam ram16s_inst_437.INIT_2 = 16'h0000;
defparam ram16s_inst_437.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_438 (
    .DO(ram16s_inst_438_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1755),
    .CLK(clk)
);

defparam ram16s_inst_438.INIT_0 = 16'h0000;
defparam ram16s_inst_438.INIT_1 = 16'h0000;
defparam ram16s_inst_438.INIT_2 = 16'h0000;
defparam ram16s_inst_438.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_439 (
    .DO(ram16s_inst_439_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1759),
    .CLK(clk)
);

defparam ram16s_inst_439.INIT_0 = 16'h0000;
defparam ram16s_inst_439.INIT_1 = 16'h0000;
defparam ram16s_inst_439.INIT_2 = 16'h0000;
defparam ram16s_inst_439.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_440 (
    .DO(ram16s_inst_440_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1763),
    .CLK(clk)
);

defparam ram16s_inst_440.INIT_0 = 16'h0000;
defparam ram16s_inst_440.INIT_1 = 16'h0000;
defparam ram16s_inst_440.INIT_2 = 16'h0000;
defparam ram16s_inst_440.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_441 (
    .DO(ram16s_inst_441_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1767),
    .CLK(clk)
);

defparam ram16s_inst_441.INIT_0 = 16'h0000;
defparam ram16s_inst_441.INIT_1 = 16'h0000;
defparam ram16s_inst_441.INIT_2 = 16'h0000;
defparam ram16s_inst_441.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_442 (
    .DO(ram16s_inst_442_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1771),
    .CLK(clk)
);

defparam ram16s_inst_442.INIT_0 = 16'h0000;
defparam ram16s_inst_442.INIT_1 = 16'h0000;
defparam ram16s_inst_442.INIT_2 = 16'h0000;
defparam ram16s_inst_442.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_443 (
    .DO(ram16s_inst_443_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1775),
    .CLK(clk)
);

defparam ram16s_inst_443.INIT_0 = 16'h0000;
defparam ram16s_inst_443.INIT_1 = 16'h0000;
defparam ram16s_inst_443.INIT_2 = 16'h0000;
defparam ram16s_inst_443.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_444 (
    .DO(ram16s_inst_444_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1779),
    .CLK(clk)
);

defparam ram16s_inst_444.INIT_0 = 16'h0000;
defparam ram16s_inst_444.INIT_1 = 16'h0000;
defparam ram16s_inst_444.INIT_2 = 16'h0000;
defparam ram16s_inst_444.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_445 (
    .DO(ram16s_inst_445_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1783),
    .CLK(clk)
);

defparam ram16s_inst_445.INIT_0 = 16'h0000;
defparam ram16s_inst_445.INIT_1 = 16'h0000;
defparam ram16s_inst_445.INIT_2 = 16'h0000;
defparam ram16s_inst_445.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_446 (
    .DO(ram16s_inst_446_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1787),
    .CLK(clk)
);

defparam ram16s_inst_446.INIT_0 = 16'h0000;
defparam ram16s_inst_446.INIT_1 = 16'h0000;
defparam ram16s_inst_446.INIT_2 = 16'h0000;
defparam ram16s_inst_446.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_447 (
    .DO(ram16s_inst_447_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1791),
    .CLK(clk)
);

defparam ram16s_inst_447.INIT_0 = 16'h0000;
defparam ram16s_inst_447.INIT_1 = 16'h0000;
defparam ram16s_inst_447.INIT_2 = 16'h0000;
defparam ram16s_inst_447.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_448 (
    .DO(ram16s_inst_448_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1795),
    .CLK(clk)
);

defparam ram16s_inst_448.INIT_0 = 16'h0000;
defparam ram16s_inst_448.INIT_1 = 16'h0000;
defparam ram16s_inst_448.INIT_2 = 16'h0000;
defparam ram16s_inst_448.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_449 (
    .DO(ram16s_inst_449_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1799),
    .CLK(clk)
);

defparam ram16s_inst_449.INIT_0 = 16'h0000;
defparam ram16s_inst_449.INIT_1 = 16'h0000;
defparam ram16s_inst_449.INIT_2 = 16'h0000;
defparam ram16s_inst_449.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_450 (
    .DO(ram16s_inst_450_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1803),
    .CLK(clk)
);

defparam ram16s_inst_450.INIT_0 = 16'h0000;
defparam ram16s_inst_450.INIT_1 = 16'h0000;
defparam ram16s_inst_450.INIT_2 = 16'h0000;
defparam ram16s_inst_450.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_451 (
    .DO(ram16s_inst_451_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1807),
    .CLK(clk)
);

defparam ram16s_inst_451.INIT_0 = 16'h0000;
defparam ram16s_inst_451.INIT_1 = 16'h0000;
defparam ram16s_inst_451.INIT_2 = 16'h0000;
defparam ram16s_inst_451.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_452 (
    .DO(ram16s_inst_452_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1811),
    .CLK(clk)
);

defparam ram16s_inst_452.INIT_0 = 16'h0000;
defparam ram16s_inst_452.INIT_1 = 16'h0000;
defparam ram16s_inst_452.INIT_2 = 16'h0000;
defparam ram16s_inst_452.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_453 (
    .DO(ram16s_inst_453_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1815),
    .CLK(clk)
);

defparam ram16s_inst_453.INIT_0 = 16'h0000;
defparam ram16s_inst_453.INIT_1 = 16'h0000;
defparam ram16s_inst_453.INIT_2 = 16'h0000;
defparam ram16s_inst_453.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_454 (
    .DO(ram16s_inst_454_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1819),
    .CLK(clk)
);

defparam ram16s_inst_454.INIT_0 = 16'h0000;
defparam ram16s_inst_454.INIT_1 = 16'h0000;
defparam ram16s_inst_454.INIT_2 = 16'h0000;
defparam ram16s_inst_454.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_455 (
    .DO(ram16s_inst_455_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1823),
    .CLK(clk)
);

defparam ram16s_inst_455.INIT_0 = 16'h0000;
defparam ram16s_inst_455.INIT_1 = 16'h0000;
defparam ram16s_inst_455.INIT_2 = 16'h0000;
defparam ram16s_inst_455.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_456 (
    .DO(ram16s_inst_456_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1827),
    .CLK(clk)
);

defparam ram16s_inst_456.INIT_0 = 16'h0000;
defparam ram16s_inst_456.INIT_1 = 16'h0000;
defparam ram16s_inst_456.INIT_2 = 16'h0000;
defparam ram16s_inst_456.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_457 (
    .DO(ram16s_inst_457_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1831),
    .CLK(clk)
);

defparam ram16s_inst_457.INIT_0 = 16'h0000;
defparam ram16s_inst_457.INIT_1 = 16'h0000;
defparam ram16s_inst_457.INIT_2 = 16'h0000;
defparam ram16s_inst_457.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_458 (
    .DO(ram16s_inst_458_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1835),
    .CLK(clk)
);

defparam ram16s_inst_458.INIT_0 = 16'h0000;
defparam ram16s_inst_458.INIT_1 = 16'h0000;
defparam ram16s_inst_458.INIT_2 = 16'h0000;
defparam ram16s_inst_458.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_459 (
    .DO(ram16s_inst_459_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1839),
    .CLK(clk)
);

defparam ram16s_inst_459.INIT_0 = 16'h0000;
defparam ram16s_inst_459.INIT_1 = 16'h0000;
defparam ram16s_inst_459.INIT_2 = 16'h0000;
defparam ram16s_inst_459.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_460 (
    .DO(ram16s_inst_460_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1843),
    .CLK(clk)
);

defparam ram16s_inst_460.INIT_0 = 16'h0000;
defparam ram16s_inst_460.INIT_1 = 16'h0000;
defparam ram16s_inst_460.INIT_2 = 16'h0000;
defparam ram16s_inst_460.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_461 (
    .DO(ram16s_inst_461_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1847),
    .CLK(clk)
);

defparam ram16s_inst_461.INIT_0 = 16'h0000;
defparam ram16s_inst_461.INIT_1 = 16'h0000;
defparam ram16s_inst_461.INIT_2 = 16'h0000;
defparam ram16s_inst_461.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_462 (
    .DO(ram16s_inst_462_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1851),
    .CLK(clk)
);

defparam ram16s_inst_462.INIT_0 = 16'h0000;
defparam ram16s_inst_462.INIT_1 = 16'h0000;
defparam ram16s_inst_462.INIT_2 = 16'h0000;
defparam ram16s_inst_462.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_463 (
    .DO(ram16s_inst_463_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1855),
    .CLK(clk)
);

defparam ram16s_inst_463.INIT_0 = 16'h0000;
defparam ram16s_inst_463.INIT_1 = 16'h0000;
defparam ram16s_inst_463.INIT_2 = 16'h0000;
defparam ram16s_inst_463.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_464 (
    .DO(ram16s_inst_464_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1859),
    .CLK(clk)
);

defparam ram16s_inst_464.INIT_0 = 16'h0000;
defparam ram16s_inst_464.INIT_1 = 16'h0000;
defparam ram16s_inst_464.INIT_2 = 16'h0000;
defparam ram16s_inst_464.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_465 (
    .DO(ram16s_inst_465_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1863),
    .CLK(clk)
);

defparam ram16s_inst_465.INIT_0 = 16'h0000;
defparam ram16s_inst_465.INIT_1 = 16'h0000;
defparam ram16s_inst_465.INIT_2 = 16'h0000;
defparam ram16s_inst_465.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_466 (
    .DO(ram16s_inst_466_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1867),
    .CLK(clk)
);

defparam ram16s_inst_466.INIT_0 = 16'h0000;
defparam ram16s_inst_466.INIT_1 = 16'h0000;
defparam ram16s_inst_466.INIT_2 = 16'h0000;
defparam ram16s_inst_466.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_467 (
    .DO(ram16s_inst_467_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1871),
    .CLK(clk)
);

defparam ram16s_inst_467.INIT_0 = 16'h0000;
defparam ram16s_inst_467.INIT_1 = 16'h0000;
defparam ram16s_inst_467.INIT_2 = 16'h0000;
defparam ram16s_inst_467.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_468 (
    .DO(ram16s_inst_468_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1875),
    .CLK(clk)
);

defparam ram16s_inst_468.INIT_0 = 16'h0000;
defparam ram16s_inst_468.INIT_1 = 16'h0000;
defparam ram16s_inst_468.INIT_2 = 16'h0000;
defparam ram16s_inst_468.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_469 (
    .DO(ram16s_inst_469_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1879),
    .CLK(clk)
);

defparam ram16s_inst_469.INIT_0 = 16'h0000;
defparam ram16s_inst_469.INIT_1 = 16'h0000;
defparam ram16s_inst_469.INIT_2 = 16'h0000;
defparam ram16s_inst_469.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_470 (
    .DO(ram16s_inst_470_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1883),
    .CLK(clk)
);

defparam ram16s_inst_470.INIT_0 = 16'h0000;
defparam ram16s_inst_470.INIT_1 = 16'h0000;
defparam ram16s_inst_470.INIT_2 = 16'h0000;
defparam ram16s_inst_470.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_471 (
    .DO(ram16s_inst_471_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1887),
    .CLK(clk)
);

defparam ram16s_inst_471.INIT_0 = 16'h000C;
defparam ram16s_inst_471.INIT_1 = 16'h0000;
defparam ram16s_inst_471.INIT_2 = 16'h0000;
defparam ram16s_inst_471.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_472 (
    .DO(ram16s_inst_472_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1891),
    .CLK(clk)
);

defparam ram16s_inst_472.INIT_0 = 16'h0000;
defparam ram16s_inst_472.INIT_1 = 16'h0000;
defparam ram16s_inst_472.INIT_2 = 16'h0000;
defparam ram16s_inst_472.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_473 (
    .DO(ram16s_inst_473_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1895),
    .CLK(clk)
);

defparam ram16s_inst_473.INIT_0 = 16'h1800;
defparam ram16s_inst_473.INIT_1 = 16'h0000;
defparam ram16s_inst_473.INIT_2 = 16'h0000;
defparam ram16s_inst_473.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_474 (
    .DO(ram16s_inst_474_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1899),
    .CLK(clk)
);

defparam ram16s_inst_474.INIT_0 = 16'h0000;
defparam ram16s_inst_474.INIT_1 = 16'h0000;
defparam ram16s_inst_474.INIT_2 = 16'h0000;
defparam ram16s_inst_474.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_475 (
    .DO(ram16s_inst_475_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1903),
    .CLK(clk)
);

defparam ram16s_inst_475.INIT_0 = 16'hFF80;
defparam ram16s_inst_475.INIT_1 = 16'h0000;
defparam ram16s_inst_475.INIT_2 = 16'h0000;
defparam ram16s_inst_475.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_476 (
    .DO(ram16s_inst_476_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1907),
    .CLK(clk)
);

defparam ram16s_inst_476.INIT_0 = 16'h000C;
defparam ram16s_inst_476.INIT_1 = 16'h0000;
defparam ram16s_inst_476.INIT_2 = 16'h0000;
defparam ram16s_inst_476.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_477 (
    .DO(ram16s_inst_477_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1911),
    .CLK(clk)
);

defparam ram16s_inst_477.INIT_0 = 16'h0000;
defparam ram16s_inst_477.INIT_1 = 16'h0000;
defparam ram16s_inst_477.INIT_2 = 16'h0000;
defparam ram16s_inst_477.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_478 (
    .DO(ram16s_inst_478_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1915),
    .CLK(clk)
);

defparam ram16s_inst_478.INIT_0 = 16'h1800;
defparam ram16s_inst_478.INIT_1 = 16'h0000;
defparam ram16s_inst_478.INIT_2 = 16'h0000;
defparam ram16s_inst_478.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_479 (
    .DO(ram16s_inst_479_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1919),
    .CLK(clk)
);

defparam ram16s_inst_479.INIT_0 = 16'h0000;
defparam ram16s_inst_479.INIT_1 = 16'h0000;
defparam ram16s_inst_479.INIT_2 = 16'h0000;
defparam ram16s_inst_479.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_480 (
    .DO(ram16s_inst_480_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1923),
    .CLK(clk)
);

defparam ram16s_inst_480.INIT_0 = 16'hFF80;
defparam ram16s_inst_480.INIT_1 = 16'h0000;
defparam ram16s_inst_480.INIT_2 = 16'h0000;
defparam ram16s_inst_480.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_481 (
    .DO(ram16s_inst_481_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1927),
    .CLK(clk)
);

defparam ram16s_inst_481.INIT_0 = 16'h000C;
defparam ram16s_inst_481.INIT_1 = 16'h0000;
defparam ram16s_inst_481.INIT_2 = 16'h0000;
defparam ram16s_inst_481.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_482 (
    .DO(ram16s_inst_482_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1931),
    .CLK(clk)
);

defparam ram16s_inst_482.INIT_0 = 16'h0000;
defparam ram16s_inst_482.INIT_1 = 16'h0000;
defparam ram16s_inst_482.INIT_2 = 16'h0000;
defparam ram16s_inst_482.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_483 (
    .DO(ram16s_inst_483_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1935),
    .CLK(clk)
);

defparam ram16s_inst_483.INIT_0 = 16'h1800;
defparam ram16s_inst_483.INIT_1 = 16'h0000;
defparam ram16s_inst_483.INIT_2 = 16'h0000;
defparam ram16s_inst_483.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_484 (
    .DO(ram16s_inst_484_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1939),
    .CLK(clk)
);

defparam ram16s_inst_484.INIT_0 = 16'h0000;
defparam ram16s_inst_484.INIT_1 = 16'h0000;
defparam ram16s_inst_484.INIT_2 = 16'h0000;
defparam ram16s_inst_484.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_485 (
    .DO(ram16s_inst_485_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1943),
    .CLK(clk)
);

defparam ram16s_inst_485.INIT_0 = 16'h1800;
defparam ram16s_inst_485.INIT_1 = 16'h0000;
defparam ram16s_inst_485.INIT_2 = 16'h0000;
defparam ram16s_inst_485.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_486 (
    .DO(ram16s_inst_486_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1947),
    .CLK(clk)
);

defparam ram16s_inst_486.INIT_0 = 16'h000C;
defparam ram16s_inst_486.INIT_1 = 16'h0000;
defparam ram16s_inst_486.INIT_2 = 16'h0000;
defparam ram16s_inst_486.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_487 (
    .DO(ram16s_inst_487_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1951),
    .CLK(clk)
);

defparam ram16s_inst_487.INIT_0 = 16'h0000;
defparam ram16s_inst_487.INIT_1 = 16'h0000;
defparam ram16s_inst_487.INIT_2 = 16'h0000;
defparam ram16s_inst_487.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_488 (
    .DO(ram16s_inst_488_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1955),
    .CLK(clk)
);

defparam ram16s_inst_488.INIT_0 = 16'h1800;
defparam ram16s_inst_488.INIT_1 = 16'h0000;
defparam ram16s_inst_488.INIT_2 = 16'h0000;
defparam ram16s_inst_488.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_489 (
    .DO(ram16s_inst_489_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1959),
    .CLK(clk)
);

defparam ram16s_inst_489.INIT_0 = 16'h0000;
defparam ram16s_inst_489.INIT_1 = 16'h0000;
defparam ram16s_inst_489.INIT_2 = 16'h0000;
defparam ram16s_inst_489.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_490 (
    .DO(ram16s_inst_490_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1963),
    .CLK(clk)
);

defparam ram16s_inst_490.INIT_0 = 16'h1800;
defparam ram16s_inst_490.INIT_1 = 16'h0000;
defparam ram16s_inst_490.INIT_2 = 16'h0000;
defparam ram16s_inst_490.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_491 (
    .DO(ram16s_inst_491_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1967),
    .CLK(clk)
);

defparam ram16s_inst_491.INIT_0 = 16'h30CC;
defparam ram16s_inst_491.INIT_1 = 16'h0000;
defparam ram16s_inst_491.INIT_2 = 16'h0000;
defparam ram16s_inst_491.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_492 (
    .DO(ram16s_inst_492_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1971),
    .CLK(clk)
);

defparam ram16s_inst_492.INIT_0 = 16'hC0E1;
defparam ram16s_inst_492.INIT_1 = 16'h0000;
defparam ram16s_inst_492.INIT_2 = 16'h0000;
defparam ram16s_inst_492.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_493 (
    .DO(ram16s_inst_493_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1975),
    .CLK(clk)
);

defparam ram16s_inst_493.INIT_0 = 16'h1981;
defparam ram16s_inst_493.INIT_1 = 16'h0000;
defparam ram16s_inst_493.INIT_2 = 16'h0000;
defparam ram16s_inst_493.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_494 (
    .DO(ram16s_inst_494_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1979),
    .CLK(clk)
);

defparam ram16s_inst_494.INIT_0 = 16'h0000;
defparam ram16s_inst_494.INIT_1 = 16'h0000;
defparam ram16s_inst_494.INIT_2 = 16'h0000;
defparam ram16s_inst_494.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_495 (
    .DO(ram16s_inst_495_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1983),
    .CLK(clk)
);

defparam ram16s_inst_495.INIT_0 = 16'h1800;
defparam ram16s_inst_495.INIT_1 = 16'h0000;
defparam ram16s_inst_495.INIT_2 = 16'h0000;
defparam ram16s_inst_495.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_496 (
    .DO(ram16s_inst_496_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1987),
    .CLK(clk)
);

defparam ram16s_inst_496.INIT_0 = 16'hF1EC;
defparam ram16s_inst_496.INIT_1 = 16'h0000;
defparam ram16s_inst_496.INIT_2 = 16'h0000;
defparam ram16s_inst_496.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_497 (
    .DO(ram16s_inst_497_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1991),
    .CLK(clk)
);

defparam ram16s_inst_497.INIT_0 = 16'hF3F9;
defparam ram16s_inst_497.INIT_1 = 16'h0000;
defparam ram16s_inst_497.INIT_2 = 16'h0000;
defparam ram16s_inst_497.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_498 (
    .DO(ram16s_inst_498_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1995),
    .CLK(clk)
);

defparam ram16s_inst_498.INIT_0 = 16'h1FC7;
defparam ram16s_inst_498.INIT_1 = 16'h0000;
defparam ram16s_inst_498.INIT_2 = 16'h0000;
defparam ram16s_inst_498.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_499 (
    .DO(ram16s_inst_499_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1999),
    .CLK(clk)
);

defparam ram16s_inst_499.INIT_0 = 16'h0000;
defparam ram16s_inst_499.INIT_1 = 16'h0000;
defparam ram16s_inst_499.INIT_2 = 16'h0000;
defparam ram16s_inst_499.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_500 (
    .DO(ram16s_inst_500_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2003),
    .CLK(clk)
);

defparam ram16s_inst_500.INIT_0 = 16'h1800;
defparam ram16s_inst_500.INIT_1 = 16'h0000;
defparam ram16s_inst_500.INIT_2 = 16'h0000;
defparam ram16s_inst_500.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_501 (
    .DO(ram16s_inst_501_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2007),
    .CLK(clk)
);

defparam ram16s_inst_501.INIT_0 = 16'h310C;
defparam ram16s_inst_501.INIT_1 = 16'h0000;
defparam ram16s_inst_501.INIT_2 = 16'h0000;
defparam ram16s_inst_501.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_502 (
    .DO(ram16s_inst_502_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2011),
    .CLK(clk)
);

defparam ram16s_inst_502.INIT_0 = 16'h0308;
defparam ram16s_inst_502.INIT_1 = 16'h0000;
defparam ram16s_inst_502.INIT_2 = 16'h0000;
defparam ram16s_inst_502.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_503 (
    .DO(ram16s_inst_503_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2015),
    .CLK(clk)
);

defparam ram16s_inst_503.INIT_0 = 16'h1866;
defparam ram16s_inst_503.INIT_1 = 16'h0000;
defparam ram16s_inst_503.INIT_2 = 16'h0000;
defparam ram16s_inst_503.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_504 (
    .DO(ram16s_inst_504_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2019),
    .CLK(clk)
);

defparam ram16s_inst_504.INIT_0 = 16'h0000;
defparam ram16s_inst_504.INIT_1 = 16'h0000;
defparam ram16s_inst_504.INIT_2 = 16'h0000;
defparam ram16s_inst_504.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_505 (
    .DO(ram16s_inst_505_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2023),
    .CLK(clk)
);

defparam ram16s_inst_505.INIT_0 = 16'h1800;
defparam ram16s_inst_505.INIT_1 = 16'h0000;
defparam ram16s_inst_505.INIT_2 = 16'h0000;
defparam ram16s_inst_505.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_506 (
    .DO(ram16s_inst_506_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2027),
    .CLK(clk)
);

defparam ram16s_inst_506.INIT_0 = 16'h330C;
defparam ram16s_inst_506.INIT_1 = 16'h0000;
defparam ram16s_inst_506.INIT_2 = 16'h0000;
defparam ram16s_inst_506.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_507 (
    .DO(ram16s_inst_507_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2031),
    .CLK(clk)
);

defparam ram16s_inst_507.INIT_0 = 16'h83FC;
defparam ram16s_inst_507.INIT_1 = 16'h0000;
defparam ram16s_inst_507.INIT_2 = 16'h0000;
defparam ram16s_inst_507.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_508 (
    .DO(ram16s_inst_508_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2035),
    .CLK(clk)
);

defparam ram16s_inst_508.INIT_0 = 16'h1867;
defparam ram16s_inst_508.INIT_1 = 16'h0000;
defparam ram16s_inst_508.INIT_2 = 16'h0000;
defparam ram16s_inst_508.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_509 (
    .DO(ram16s_inst_509_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2039),
    .CLK(clk)
);

defparam ram16s_inst_509.INIT_0 = 16'h0000;
defparam ram16s_inst_509.INIT_1 = 16'h0000;
defparam ram16s_inst_509.INIT_2 = 16'h0000;
defparam ram16s_inst_509.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_510 (
    .DO(ram16s_inst_510_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2043),
    .CLK(clk)
);

defparam ram16s_inst_510.INIT_0 = 16'h1800;
defparam ram16s_inst_510.INIT_1 = 16'h0000;
defparam ram16s_inst_510.INIT_2 = 16'h0000;
defparam ram16s_inst_510.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_511 (
    .DO(ram16s_inst_511_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2047),
    .CLK(clk)
);

defparam ram16s_inst_511.INIT_0 = 16'h330C;
defparam ram16s_inst_511.INIT_1 = 16'h0000;
defparam ram16s_inst_511.INIT_2 = 16'h0000;
defparam ram16s_inst_511.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_512 (
    .DO(ram16s_inst_512_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2051),
    .CLK(clk)
);

defparam ram16s_inst_512.INIT_0 = 16'h100C;
defparam ram16s_inst_512.INIT_1 = 16'h0000;
defparam ram16s_inst_512.INIT_2 = 16'h0000;
defparam ram16s_inst_512.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_513 (
    .DO(ram16s_inst_513_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2055),
    .CLK(clk)
);

defparam ram16s_inst_513.INIT_0 = 16'h1826;
defparam ram16s_inst_513.INIT_1 = 16'h0000;
defparam ram16s_inst_513.INIT_2 = 16'h0000;
defparam ram16s_inst_513.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_514 (
    .DO(ram16s_inst_514_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2059),
    .CLK(clk)
);

defparam ram16s_inst_514.INIT_0 = 16'h0000;
defparam ram16s_inst_514.INIT_1 = 16'h0000;
defparam ram16s_inst_514.INIT_2 = 16'h0000;
defparam ram16s_inst_514.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_515 (
    .DO(ram16s_inst_515_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2063),
    .CLK(clk)
);

defparam ram16s_inst_515.INIT_0 = 16'h1800;
defparam ram16s_inst_515.INIT_1 = 16'h0000;
defparam ram16s_inst_515.INIT_2 = 16'h0000;
defparam ram16s_inst_515.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_516 (
    .DO(ram16s_inst_516_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2067),
    .CLK(clk)
);

defparam ram16s_inst_516.INIT_0 = 16'h330C;
defparam ram16s_inst_516.INIT_1 = 16'h0000;
defparam ram16s_inst_516.INIT_2 = 16'h0000;
defparam ram16s_inst_516.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_517 (
    .DO(ram16s_inst_517_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2071),
    .CLK(clk)
);

defparam ram16s_inst_517.INIT_0 = 16'h1018;
defparam ram16s_inst_517.INIT_1 = 16'h0000;
defparam ram16s_inst_517.INIT_2 = 16'h0000;
defparam ram16s_inst_517.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_518 (
    .DO(ram16s_inst_518_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2075),
    .CLK(clk)
);

defparam ram16s_inst_518.INIT_0 = 16'h1866;
defparam ram16s_inst_518.INIT_1 = 16'h0000;
defparam ram16s_inst_518.INIT_2 = 16'h0000;
defparam ram16s_inst_518.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_519 (
    .DO(ram16s_inst_519_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2079),
    .CLK(clk)
);

defparam ram16s_inst_519.INIT_0 = 16'h0000;
defparam ram16s_inst_519.INIT_1 = 16'h0000;
defparam ram16s_inst_519.INIT_2 = 16'h0000;
defparam ram16s_inst_519.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_520 (
    .DO(ram16s_inst_520_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2083),
    .CLK(clk)
);

defparam ram16s_inst_520.INIT_0 = 16'h1800;
defparam ram16s_inst_520.INIT_1 = 16'h0000;
defparam ram16s_inst_520.INIT_2 = 16'h0000;
defparam ram16s_inst_520.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_521 (
    .DO(ram16s_inst_521_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2087),
    .CLK(clk)
);

defparam ram16s_inst_521.INIT_0 = 16'h330C;
defparam ram16s_inst_521.INIT_1 = 16'h0000;
defparam ram16s_inst_521.INIT_2 = 16'h0000;
defparam ram16s_inst_521.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_522 (
    .DO(ram16s_inst_522_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2091),
    .CLK(clk)
);

defparam ram16s_inst_522.INIT_0 = 16'hF3F8;
defparam ram16s_inst_522.INIT_1 = 16'h0000;
defparam ram16s_inst_522.INIT_2 = 16'h0000;
defparam ram16s_inst_522.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_523 (
    .DO(ram16s_inst_523_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2095),
    .CLK(clk)
);

defparam ram16s_inst_523.INIT_0 = 16'h1FE6;
defparam ram16s_inst_523.INIT_1 = 16'h0000;
defparam ram16s_inst_523.INIT_2 = 16'h0000;
defparam ram16s_inst_523.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_524 (
    .DO(ram16s_inst_524_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2099),
    .CLK(clk)
);

defparam ram16s_inst_524.INIT_0 = 16'h0000;
defparam ram16s_inst_524.INIT_1 = 16'h0000;
defparam ram16s_inst_524.INIT_2 = 16'h0000;
defparam ram16s_inst_524.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_525 (
    .DO(ram16s_inst_525_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2103),
    .CLK(clk)
);

defparam ram16s_inst_525.INIT_0 = 16'h1800;
defparam ram16s_inst_525.INIT_1 = 16'h0000;
defparam ram16s_inst_525.INIT_2 = 16'h0000;
defparam ram16s_inst_525.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_526 (
    .DO(ram16s_inst_526_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2107),
    .CLK(clk)
);

defparam ram16s_inst_526.INIT_0 = 16'h330C;
defparam ram16s_inst_526.INIT_1 = 16'h0000;
defparam ram16s_inst_526.INIT_2 = 16'h0000;
defparam ram16s_inst_526.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_527 (
    .DO(ram16s_inst_527_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2111),
    .CLK(clk)
);

defparam ram16s_inst_527.INIT_0 = 16'h60E0;
defparam ram16s_inst_527.INIT_1 = 16'h0000;
defparam ram16s_inst_527.INIT_2 = 16'h0000;
defparam ram16s_inst_527.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_528 (
    .DO(ram16s_inst_528_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2115),
    .CLK(clk)
);

defparam ram16s_inst_528.INIT_0 = 16'h1986;
defparam ram16s_inst_528.INIT_1 = 16'h0000;
defparam ram16s_inst_528.INIT_2 = 16'h0000;
defparam ram16s_inst_528.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_529 (
    .DO(ram16s_inst_529_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2119),
    .CLK(clk)
);

defparam ram16s_inst_529.INIT_0 = 16'h0000;
defparam ram16s_inst_529.INIT_1 = 16'h0000;
defparam ram16s_inst_529.INIT_2 = 16'h0000;
defparam ram16s_inst_529.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_530 (
    .DO(ram16s_inst_530_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2123),
    .CLK(clk)
);

defparam ram16s_inst_530.INIT_0 = 16'h0000;
defparam ram16s_inst_530.INIT_1 = 16'h0000;
defparam ram16s_inst_530.INIT_2 = 16'h0000;
defparam ram16s_inst_530.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_531 (
    .DO(ram16s_inst_531_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2127),
    .CLK(clk)
);

defparam ram16s_inst_531.INIT_0 = 16'h0000;
defparam ram16s_inst_531.INIT_1 = 16'h0000;
defparam ram16s_inst_531.INIT_2 = 16'h0000;
defparam ram16s_inst_531.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_532 (
    .DO(ram16s_inst_532_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2131),
    .CLK(clk)
);

defparam ram16s_inst_532.INIT_0 = 16'h0000;
defparam ram16s_inst_532.INIT_1 = 16'h0000;
defparam ram16s_inst_532.INIT_2 = 16'h0000;
defparam ram16s_inst_532.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_533 (
    .DO(ram16s_inst_533_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2135),
    .CLK(clk)
);

defparam ram16s_inst_533.INIT_0 = 16'h0000;
defparam ram16s_inst_533.INIT_1 = 16'h0000;
defparam ram16s_inst_533.INIT_2 = 16'h0000;
defparam ram16s_inst_533.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_534 (
    .DO(ram16s_inst_534_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2139),
    .CLK(clk)
);

defparam ram16s_inst_534.INIT_0 = 16'h0000;
defparam ram16s_inst_534.INIT_1 = 16'h0000;
defparam ram16s_inst_534.INIT_2 = 16'h0000;
defparam ram16s_inst_534.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_535 (
    .DO(ram16s_inst_535_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2143),
    .CLK(clk)
);

defparam ram16s_inst_535.INIT_0 = 16'h0000;
defparam ram16s_inst_535.INIT_1 = 16'h0000;
defparam ram16s_inst_535.INIT_2 = 16'h0000;
defparam ram16s_inst_535.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_536 (
    .DO(ram16s_inst_536_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2147),
    .CLK(clk)
);

defparam ram16s_inst_536.INIT_0 = 16'h0000;
defparam ram16s_inst_536.INIT_1 = 16'h0000;
defparam ram16s_inst_536.INIT_2 = 16'h0000;
defparam ram16s_inst_536.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_537 (
    .DO(ram16s_inst_537_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2151),
    .CLK(clk)
);

defparam ram16s_inst_537.INIT_0 = 16'h0000;
defparam ram16s_inst_537.INIT_1 = 16'h0000;
defparam ram16s_inst_537.INIT_2 = 16'h0000;
defparam ram16s_inst_537.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_538 (
    .DO(ram16s_inst_538_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2155),
    .CLK(clk)
);

defparam ram16s_inst_538.INIT_0 = 16'h0000;
defparam ram16s_inst_538.INIT_1 = 16'h0000;
defparam ram16s_inst_538.INIT_2 = 16'h0000;
defparam ram16s_inst_538.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_539 (
    .DO(ram16s_inst_539_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2159),
    .CLK(clk)
);

defparam ram16s_inst_539.INIT_0 = 16'h0000;
defparam ram16s_inst_539.INIT_1 = 16'h0000;
defparam ram16s_inst_539.INIT_2 = 16'h0000;
defparam ram16s_inst_539.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_540 (
    .DO(ram16s_inst_540_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2163),
    .CLK(clk)
);

defparam ram16s_inst_540.INIT_0 = 16'h0000;
defparam ram16s_inst_540.INIT_1 = 16'h0000;
defparam ram16s_inst_540.INIT_2 = 16'h0000;
defparam ram16s_inst_540.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_541 (
    .DO(ram16s_inst_541_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2167),
    .CLK(clk)
);

defparam ram16s_inst_541.INIT_0 = 16'h0000;
defparam ram16s_inst_541.INIT_1 = 16'h0000;
defparam ram16s_inst_541.INIT_2 = 16'h0000;
defparam ram16s_inst_541.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_542 (
    .DO(ram16s_inst_542_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2171),
    .CLK(clk)
);

defparam ram16s_inst_542.INIT_0 = 16'h0000;
defparam ram16s_inst_542.INIT_1 = 16'h0000;
defparam ram16s_inst_542.INIT_2 = 16'h0000;
defparam ram16s_inst_542.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_543 (
    .DO(ram16s_inst_543_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2175),
    .CLK(clk)
);

defparam ram16s_inst_543.INIT_0 = 16'h0000;
defparam ram16s_inst_543.INIT_1 = 16'h0000;
defparam ram16s_inst_543.INIT_2 = 16'h0000;
defparam ram16s_inst_543.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_544 (
    .DO(ram16s_inst_544_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2179),
    .CLK(clk)
);

defparam ram16s_inst_544.INIT_0 = 16'h0000;
defparam ram16s_inst_544.INIT_1 = 16'h0000;
defparam ram16s_inst_544.INIT_2 = 16'h0000;
defparam ram16s_inst_544.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_545 (
    .DO(ram16s_inst_545_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2183),
    .CLK(clk)
);

defparam ram16s_inst_545.INIT_0 = 16'h0000;
defparam ram16s_inst_545.INIT_1 = 16'h0000;
defparam ram16s_inst_545.INIT_2 = 16'h0000;
defparam ram16s_inst_545.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_546 (
    .DO(ram16s_inst_546_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2187),
    .CLK(clk)
);

defparam ram16s_inst_546.INIT_0 = 16'h0000;
defparam ram16s_inst_546.INIT_1 = 16'h0000;
defparam ram16s_inst_546.INIT_2 = 16'h0000;
defparam ram16s_inst_546.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_547 (
    .DO(ram16s_inst_547_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2191),
    .CLK(clk)
);

defparam ram16s_inst_547.INIT_0 = 16'h0000;
defparam ram16s_inst_547.INIT_1 = 16'h0000;
defparam ram16s_inst_547.INIT_2 = 16'h0000;
defparam ram16s_inst_547.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_548 (
    .DO(ram16s_inst_548_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2195),
    .CLK(clk)
);

defparam ram16s_inst_548.INIT_0 = 16'h0000;
defparam ram16s_inst_548.INIT_1 = 16'h0000;
defparam ram16s_inst_548.INIT_2 = 16'h0000;
defparam ram16s_inst_548.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_549 (
    .DO(ram16s_inst_549_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2199),
    .CLK(clk)
);

defparam ram16s_inst_549.INIT_0 = 16'h0000;
defparam ram16s_inst_549.INIT_1 = 16'h0000;
defparam ram16s_inst_549.INIT_2 = 16'h0000;
defparam ram16s_inst_549.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_550 (
    .DO(ram16s_inst_550_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2203),
    .CLK(clk)
);

defparam ram16s_inst_550.INIT_0 = 16'h0000;
defparam ram16s_inst_550.INIT_1 = 16'h0000;
defparam ram16s_inst_550.INIT_2 = 16'h0000;
defparam ram16s_inst_550.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_551 (
    .DO(ram16s_inst_551_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2207),
    .CLK(clk)
);

defparam ram16s_inst_551.INIT_0 = 16'h0000;
defparam ram16s_inst_551.INIT_1 = 16'h0000;
defparam ram16s_inst_551.INIT_2 = 16'h0000;
defparam ram16s_inst_551.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_552 (
    .DO(ram16s_inst_552_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2211),
    .CLK(clk)
);

defparam ram16s_inst_552.INIT_0 = 16'h0000;
defparam ram16s_inst_552.INIT_1 = 16'h0000;
defparam ram16s_inst_552.INIT_2 = 16'h0000;
defparam ram16s_inst_552.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_553 (
    .DO(ram16s_inst_553_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2215),
    .CLK(clk)
);

defparam ram16s_inst_553.INIT_0 = 16'h0000;
defparam ram16s_inst_553.INIT_1 = 16'h0000;
defparam ram16s_inst_553.INIT_2 = 16'h0000;
defparam ram16s_inst_553.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_554 (
    .DO(ram16s_inst_554_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2219),
    .CLK(clk)
);

defparam ram16s_inst_554.INIT_0 = 16'h0000;
defparam ram16s_inst_554.INIT_1 = 16'h0000;
defparam ram16s_inst_554.INIT_2 = 16'h0000;
defparam ram16s_inst_554.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_555 (
    .DO(ram16s_inst_555_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2223),
    .CLK(clk)
);

defparam ram16s_inst_555.INIT_0 = 16'h0000;
defparam ram16s_inst_555.INIT_1 = 16'h0000;
defparam ram16s_inst_555.INIT_2 = 16'h0000;
defparam ram16s_inst_555.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_556 (
    .DO(ram16s_inst_556_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2227),
    .CLK(clk)
);

defparam ram16s_inst_556.INIT_0 = 16'h0000;
defparam ram16s_inst_556.INIT_1 = 16'h0000;
defparam ram16s_inst_556.INIT_2 = 16'h0000;
defparam ram16s_inst_556.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_557 (
    .DO(ram16s_inst_557_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2231),
    .CLK(clk)
);

defparam ram16s_inst_557.INIT_0 = 16'h0000;
defparam ram16s_inst_557.INIT_1 = 16'h0000;
defparam ram16s_inst_557.INIT_2 = 16'h0000;
defparam ram16s_inst_557.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_558 (
    .DO(ram16s_inst_558_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2235),
    .CLK(clk)
);

defparam ram16s_inst_558.INIT_0 = 16'h0000;
defparam ram16s_inst_558.INIT_1 = 16'h0000;
defparam ram16s_inst_558.INIT_2 = 16'h0000;
defparam ram16s_inst_558.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_559 (
    .DO(ram16s_inst_559_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2239),
    .CLK(clk)
);

defparam ram16s_inst_559.INIT_0 = 16'h0000;
defparam ram16s_inst_559.INIT_1 = 16'h0000;
defparam ram16s_inst_559.INIT_2 = 16'h0000;
defparam ram16s_inst_559.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_560 (
    .DO(ram16s_inst_560_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2243),
    .CLK(clk)
);

defparam ram16s_inst_560.INIT_0 = 16'h0000;
defparam ram16s_inst_560.INIT_1 = 16'h0000;
defparam ram16s_inst_560.INIT_2 = 16'h0000;
defparam ram16s_inst_560.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_561 (
    .DO(ram16s_inst_561_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2247),
    .CLK(clk)
);

defparam ram16s_inst_561.INIT_0 = 16'h0000;
defparam ram16s_inst_561.INIT_1 = 16'h0000;
defparam ram16s_inst_561.INIT_2 = 16'h0000;
defparam ram16s_inst_561.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_562 (
    .DO(ram16s_inst_562_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2251),
    .CLK(clk)
);

defparam ram16s_inst_562.INIT_0 = 16'h0000;
defparam ram16s_inst_562.INIT_1 = 16'h0000;
defparam ram16s_inst_562.INIT_2 = 16'h0000;
defparam ram16s_inst_562.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_563 (
    .DO(ram16s_inst_563_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2255),
    .CLK(clk)
);

defparam ram16s_inst_563.INIT_0 = 16'h0000;
defparam ram16s_inst_563.INIT_1 = 16'h0000;
defparam ram16s_inst_563.INIT_2 = 16'h0000;
defparam ram16s_inst_563.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_564 (
    .DO(ram16s_inst_564_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2259),
    .CLK(clk)
);

defparam ram16s_inst_564.INIT_0 = 16'h0000;
defparam ram16s_inst_564.INIT_1 = 16'h0000;
defparam ram16s_inst_564.INIT_2 = 16'h0000;
defparam ram16s_inst_564.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_565 (
    .DO(ram16s_inst_565_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2263),
    .CLK(clk)
);

defparam ram16s_inst_565.INIT_0 = 16'h0000;
defparam ram16s_inst_565.INIT_1 = 16'h0000;
defparam ram16s_inst_565.INIT_2 = 16'hFE00;
defparam ram16s_inst_565.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_566 (
    .DO(ram16s_inst_566_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2267),
    .CLK(clk)
);

defparam ram16s_inst_566.INIT_0 = 16'h0000;
defparam ram16s_inst_566.INIT_1 = 16'h0000;
defparam ram16s_inst_566.INIT_2 = 16'h87F0;
defparam ram16s_inst_566.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_567 (
    .DO(ram16s_inst_567_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2271),
    .CLK(clk)
);

defparam ram16s_inst_567.INIT_0 = 16'h0000;
defparam ram16s_inst_567.INIT_1 = 16'h0000;
defparam ram16s_inst_567.INIT_2 = 16'hFC3F;
defparam ram16s_inst_567.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_568 (
    .DO(ram16s_inst_568_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2275),
    .CLK(clk)
);

defparam ram16s_inst_568.INIT_0 = 16'h0000;
defparam ram16s_inst_568.INIT_1 = 16'h0000;
defparam ram16s_inst_568.INIT_2 = 16'h0001;
defparam ram16s_inst_568.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_569 (
    .DO(ram16s_inst_569_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2279),
    .CLK(clk)
);

defparam ram16s_inst_569.INIT_0 = 16'h0000;
defparam ram16s_inst_569.INIT_1 = 16'h0000;
defparam ram16s_inst_569.INIT_2 = 16'h0000;
defparam ram16s_inst_569.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_570 (
    .DO(ram16s_inst_570_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2283),
    .CLK(clk)
);

defparam ram16s_inst_570.INIT_0 = 16'h0000;
defparam ram16s_inst_570.INIT_1 = 16'h0000;
defparam ram16s_inst_570.INIT_2 = 16'hFE00;
defparam ram16s_inst_570.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_571 (
    .DO(ram16s_inst_571_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2287),
    .CLK(clk)
);

defparam ram16s_inst_571.INIT_0 = 16'h0000;
defparam ram16s_inst_571.INIT_1 = 16'h0000;
defparam ram16s_inst_571.INIT_2 = 16'h87F0;
defparam ram16s_inst_571.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_572 (
    .DO(ram16s_inst_572_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2291),
    .CLK(clk)
);

defparam ram16s_inst_572.INIT_0 = 16'h0000;
defparam ram16s_inst_572.INIT_1 = 16'h0000;
defparam ram16s_inst_572.INIT_2 = 16'hFC3F;
defparam ram16s_inst_572.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_573 (
    .DO(ram16s_inst_573_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2295),
    .CLK(clk)
);

defparam ram16s_inst_573.INIT_0 = 16'h0000;
defparam ram16s_inst_573.INIT_1 = 16'h0000;
defparam ram16s_inst_573.INIT_2 = 16'h0001;
defparam ram16s_inst_573.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_574 (
    .DO(ram16s_inst_574_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2299),
    .CLK(clk)
);

defparam ram16s_inst_574.INIT_0 = 16'h0000;
defparam ram16s_inst_574.INIT_1 = 16'h0000;
defparam ram16s_inst_574.INIT_2 = 16'h0000;
defparam ram16s_inst_574.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_575 (
    .DO(ram16s_inst_575_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2303),
    .CLK(clk)
);

defparam ram16s_inst_575.INIT_0 = 16'h0000;
defparam ram16s_inst_575.INIT_1 = 16'h0000;
defparam ram16s_inst_575.INIT_2 = 16'hFE00;
defparam ram16s_inst_575.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_576 (
    .DO(ram16s_inst_576_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2307),
    .CLK(clk)
);

defparam ram16s_inst_576.INIT_0 = 16'h0000;
defparam ram16s_inst_576.INIT_1 = 16'h0000;
defparam ram16s_inst_576.INIT_2 = 16'h87F0;
defparam ram16s_inst_576.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_577 (
    .DO(ram16s_inst_577_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2311),
    .CLK(clk)
);

defparam ram16s_inst_577.INIT_0 = 16'h0000;
defparam ram16s_inst_577.INIT_1 = 16'h0000;
defparam ram16s_inst_577.INIT_2 = 16'hFC3F;
defparam ram16s_inst_577.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_578 (
    .DO(ram16s_inst_578_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2315),
    .CLK(clk)
);

defparam ram16s_inst_578.INIT_0 = 16'h0000;
defparam ram16s_inst_578.INIT_1 = 16'h0000;
defparam ram16s_inst_578.INIT_2 = 16'h0001;
defparam ram16s_inst_578.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_579 (
    .DO(ram16s_inst_579_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2319),
    .CLK(clk)
);

defparam ram16s_inst_579.INIT_0 = 16'h0000;
defparam ram16s_inst_579.INIT_1 = 16'h0000;
defparam ram16s_inst_579.INIT_2 = 16'h0000;
defparam ram16s_inst_579.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_580 (
    .DO(ram16s_inst_580_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2323),
    .CLK(clk)
);

defparam ram16s_inst_580.INIT_0 = 16'h0000;
defparam ram16s_inst_580.INIT_1 = 16'h0000;
defparam ram16s_inst_580.INIT_2 = 16'hFE00;
defparam ram16s_inst_580.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_581 (
    .DO(ram16s_inst_581_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2327),
    .CLK(clk)
);

defparam ram16s_inst_581.INIT_0 = 16'h0000;
defparam ram16s_inst_581.INIT_1 = 16'h0000;
defparam ram16s_inst_581.INIT_2 = 16'h87F0;
defparam ram16s_inst_581.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_582 (
    .DO(ram16s_inst_582_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2331),
    .CLK(clk)
);

defparam ram16s_inst_582.INIT_0 = 16'h0000;
defparam ram16s_inst_582.INIT_1 = 16'h0000;
defparam ram16s_inst_582.INIT_2 = 16'hFC3F;
defparam ram16s_inst_582.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_583 (
    .DO(ram16s_inst_583_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2335),
    .CLK(clk)
);

defparam ram16s_inst_583.INIT_0 = 16'h0000;
defparam ram16s_inst_583.INIT_1 = 16'h0000;
defparam ram16s_inst_583.INIT_2 = 16'h0001;
defparam ram16s_inst_583.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_584 (
    .DO(ram16s_inst_584_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2339),
    .CLK(clk)
);

defparam ram16s_inst_584.INIT_0 = 16'h0000;
defparam ram16s_inst_584.INIT_1 = 16'h0000;
defparam ram16s_inst_584.INIT_2 = 16'h0000;
defparam ram16s_inst_584.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_585 (
    .DO(ram16s_inst_585_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2343),
    .CLK(clk)
);

defparam ram16s_inst_585.INIT_0 = 16'h0000;
defparam ram16s_inst_585.INIT_1 = 16'h0000;
defparam ram16s_inst_585.INIT_2 = 16'hFE00;
defparam ram16s_inst_585.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_586 (
    .DO(ram16s_inst_586_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2347),
    .CLK(clk)
);

defparam ram16s_inst_586.INIT_0 = 16'h0000;
defparam ram16s_inst_586.INIT_1 = 16'h0000;
defparam ram16s_inst_586.INIT_2 = 16'h87F0;
defparam ram16s_inst_586.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_587 (
    .DO(ram16s_inst_587_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2351),
    .CLK(clk)
);

defparam ram16s_inst_587.INIT_0 = 16'h0000;
defparam ram16s_inst_587.INIT_1 = 16'h0000;
defparam ram16s_inst_587.INIT_2 = 16'hFC3F;
defparam ram16s_inst_587.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_588 (
    .DO(ram16s_inst_588_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2355),
    .CLK(clk)
);

defparam ram16s_inst_588.INIT_0 = 16'h0000;
defparam ram16s_inst_588.INIT_1 = 16'h0000;
defparam ram16s_inst_588.INIT_2 = 16'h0001;
defparam ram16s_inst_588.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_589 (
    .DO(ram16s_inst_589_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2359),
    .CLK(clk)
);

defparam ram16s_inst_589.INIT_0 = 16'h0000;
defparam ram16s_inst_589.INIT_1 = 16'h0000;
defparam ram16s_inst_589.INIT_2 = 16'h0000;
defparam ram16s_inst_589.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_590 (
    .DO(ram16s_inst_590_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2363),
    .CLK(clk)
);

defparam ram16s_inst_590.INIT_0 = 16'h0000;
defparam ram16s_inst_590.INIT_1 = 16'h0000;
defparam ram16s_inst_590.INIT_2 = 16'hFE00;
defparam ram16s_inst_590.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_591 (
    .DO(ram16s_inst_591_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2367),
    .CLK(clk)
);

defparam ram16s_inst_591.INIT_0 = 16'h0000;
defparam ram16s_inst_591.INIT_1 = 16'h0000;
defparam ram16s_inst_591.INIT_2 = 16'h87F0;
defparam ram16s_inst_591.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_592 (
    .DO(ram16s_inst_592_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2371),
    .CLK(clk)
);

defparam ram16s_inst_592.INIT_0 = 16'h0000;
defparam ram16s_inst_592.INIT_1 = 16'h0000;
defparam ram16s_inst_592.INIT_2 = 16'hFC3F;
defparam ram16s_inst_592.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_593 (
    .DO(ram16s_inst_593_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2375),
    .CLK(clk)
);

defparam ram16s_inst_593.INIT_0 = 16'h0000;
defparam ram16s_inst_593.INIT_1 = 16'h0000;
defparam ram16s_inst_593.INIT_2 = 16'h0001;
defparam ram16s_inst_593.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_594 (
    .DO(ram16s_inst_594_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2379),
    .CLK(clk)
);

defparam ram16s_inst_594.INIT_0 = 16'h0000;
defparam ram16s_inst_594.INIT_1 = 16'h0000;
defparam ram16s_inst_594.INIT_2 = 16'h0000;
defparam ram16s_inst_594.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_595 (
    .DO(ram16s_inst_595_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2383),
    .CLK(clk)
);

defparam ram16s_inst_595.INIT_0 = 16'h0000;
defparam ram16s_inst_595.INIT_1 = 16'h0000;
defparam ram16s_inst_595.INIT_2 = 16'h0000;
defparam ram16s_inst_595.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_596 (
    .DO(ram16s_inst_596_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2387),
    .CLK(clk)
);

defparam ram16s_inst_596.INIT_0 = 16'h0000;
defparam ram16s_inst_596.INIT_1 = 16'h0000;
defparam ram16s_inst_596.INIT_2 = 16'h0000;
defparam ram16s_inst_596.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_597 (
    .DO(ram16s_inst_597_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2391),
    .CLK(clk)
);

defparam ram16s_inst_597.INIT_0 = 16'h0000;
defparam ram16s_inst_597.INIT_1 = 16'h0000;
defparam ram16s_inst_597.INIT_2 = 16'h0000;
defparam ram16s_inst_597.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_598 (
    .DO(ram16s_inst_598_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2395),
    .CLK(clk)
);

defparam ram16s_inst_598.INIT_0 = 16'h0000;
defparam ram16s_inst_598.INIT_1 = 16'h0000;
defparam ram16s_inst_598.INIT_2 = 16'h0000;
defparam ram16s_inst_598.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_599 (
    .DO(ram16s_inst_599_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2399),
    .CLK(clk)
);

defparam ram16s_inst_599.INIT_0 = 16'h0000;
defparam ram16s_inst_599.INIT_1 = 16'h0000;
defparam ram16s_inst_599.INIT_2 = 16'h0000;
defparam ram16s_inst_599.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_600 (
    .DO(ram16s_inst_600_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2403),
    .CLK(clk)
);

defparam ram16s_inst_600.INIT_0 = 16'h0000;
defparam ram16s_inst_600.INIT_1 = 16'h0000;
defparam ram16s_inst_600.INIT_2 = 16'h0000;
defparam ram16s_inst_600.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_601 (
    .DO(ram16s_inst_601_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2407),
    .CLK(clk)
);

defparam ram16s_inst_601.INIT_0 = 16'h0000;
defparam ram16s_inst_601.INIT_1 = 16'h0000;
defparam ram16s_inst_601.INIT_2 = 16'h0000;
defparam ram16s_inst_601.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_602 (
    .DO(ram16s_inst_602_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2411),
    .CLK(clk)
);

defparam ram16s_inst_602.INIT_0 = 16'h0000;
defparam ram16s_inst_602.INIT_1 = 16'h0000;
defparam ram16s_inst_602.INIT_2 = 16'h0000;
defparam ram16s_inst_602.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_603 (
    .DO(ram16s_inst_603_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2415),
    .CLK(clk)
);

defparam ram16s_inst_603.INIT_0 = 16'h0000;
defparam ram16s_inst_603.INIT_1 = 16'h0000;
defparam ram16s_inst_603.INIT_2 = 16'h0000;
defparam ram16s_inst_603.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_604 (
    .DO(ram16s_inst_604_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2419),
    .CLK(clk)
);

defparam ram16s_inst_604.INIT_0 = 16'h0000;
defparam ram16s_inst_604.INIT_1 = 16'h0000;
defparam ram16s_inst_604.INIT_2 = 16'h0000;
defparam ram16s_inst_604.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_605 (
    .DO(ram16s_inst_605_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2423),
    .CLK(clk)
);

defparam ram16s_inst_605.INIT_0 = 16'h0000;
defparam ram16s_inst_605.INIT_1 = 16'h0000;
defparam ram16s_inst_605.INIT_2 = 16'h0000;
defparam ram16s_inst_605.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_606 (
    .DO(ram16s_inst_606_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2427),
    .CLK(clk)
);

defparam ram16s_inst_606.INIT_0 = 16'h0000;
defparam ram16s_inst_606.INIT_1 = 16'h0000;
defparam ram16s_inst_606.INIT_2 = 16'h0000;
defparam ram16s_inst_606.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_607 (
    .DO(ram16s_inst_607_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2431),
    .CLK(clk)
);

defparam ram16s_inst_607.INIT_0 = 16'h0000;
defparam ram16s_inst_607.INIT_1 = 16'h0000;
defparam ram16s_inst_607.INIT_2 = 16'h0000;
defparam ram16s_inst_607.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_608 (
    .DO(ram16s_inst_608_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2435),
    .CLK(clk)
);

defparam ram16s_inst_608.INIT_0 = 16'h0000;
defparam ram16s_inst_608.INIT_1 = 16'h0000;
defparam ram16s_inst_608.INIT_2 = 16'h0000;
defparam ram16s_inst_608.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_609 (
    .DO(ram16s_inst_609_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2439),
    .CLK(clk)
);

defparam ram16s_inst_609.INIT_0 = 16'h0000;
defparam ram16s_inst_609.INIT_1 = 16'h0000;
defparam ram16s_inst_609.INIT_2 = 16'h0000;
defparam ram16s_inst_609.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_610 (
    .DO(ram16s_inst_610_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2443),
    .CLK(clk)
);

defparam ram16s_inst_610.INIT_0 = 16'h0000;
defparam ram16s_inst_610.INIT_1 = 16'h0000;
defparam ram16s_inst_610.INIT_2 = 16'h0000;
defparam ram16s_inst_610.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_611 (
    .DO(ram16s_inst_611_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2447),
    .CLK(clk)
);

defparam ram16s_inst_611.INIT_0 = 16'h0000;
defparam ram16s_inst_611.INIT_1 = 16'h0000;
defparam ram16s_inst_611.INIT_2 = 16'h0000;
defparam ram16s_inst_611.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_612 (
    .DO(ram16s_inst_612_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2451),
    .CLK(clk)
);

defparam ram16s_inst_612.INIT_0 = 16'h0000;
defparam ram16s_inst_612.INIT_1 = 16'h0000;
defparam ram16s_inst_612.INIT_2 = 16'h0000;
defparam ram16s_inst_612.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_613 (
    .DO(ram16s_inst_613_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2455),
    .CLK(clk)
);

defparam ram16s_inst_613.INIT_0 = 16'h0000;
defparam ram16s_inst_613.INIT_1 = 16'h0000;
defparam ram16s_inst_613.INIT_2 = 16'h0000;
defparam ram16s_inst_613.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_614 (
    .DO(ram16s_inst_614_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2459),
    .CLK(clk)
);

defparam ram16s_inst_614.INIT_0 = 16'h0000;
defparam ram16s_inst_614.INIT_1 = 16'h0000;
defparam ram16s_inst_614.INIT_2 = 16'h0000;
defparam ram16s_inst_614.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_615 (
    .DO(ram16s_inst_615_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2463),
    .CLK(clk)
);

defparam ram16s_inst_615.INIT_0 = 16'h0000;
defparam ram16s_inst_615.INIT_1 = 16'h0000;
defparam ram16s_inst_615.INIT_2 = 16'hFE00;
defparam ram16s_inst_615.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_616 (
    .DO(ram16s_inst_616_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2467),
    .CLK(clk)
);

defparam ram16s_inst_616.INIT_0 = 16'h0000;
defparam ram16s_inst_616.INIT_1 = 16'h8000;
defparam ram16s_inst_616.INIT_2 = 16'h07F0;
defparam ram16s_inst_616.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_617 (
    .DO(ram16s_inst_617_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2471),
    .CLK(clk)
);

defparam ram16s_inst_617.INIT_0 = 16'h0000;
defparam ram16s_inst_617.INIT_1 = 16'hFC3F;
defparam ram16s_inst_617.INIT_2 = 16'h0000;
defparam ram16s_inst_617.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_618 (
    .DO(ram16s_inst_618_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2475),
    .CLK(clk)
);

defparam ram16s_inst_618.INIT_0 = 16'h0000;
defparam ram16s_inst_618.INIT_1 = 16'h0001;
defparam ram16s_inst_618.INIT_2 = 16'h0000;
defparam ram16s_inst_618.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_619 (
    .DO(ram16s_inst_619_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2479),
    .CLK(clk)
);

defparam ram16s_inst_619.INIT_0 = 16'h0000;
defparam ram16s_inst_619.INIT_1 = 16'h0000;
defparam ram16s_inst_619.INIT_2 = 16'h0000;
defparam ram16s_inst_619.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_620 (
    .DO(ram16s_inst_620_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2483),
    .CLK(clk)
);

defparam ram16s_inst_620.INIT_0 = 16'h0000;
defparam ram16s_inst_620.INIT_1 = 16'h0000;
defparam ram16s_inst_620.INIT_2 = 16'hFE00;
defparam ram16s_inst_620.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_621 (
    .DO(ram16s_inst_621_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2487),
    .CLK(clk)
);

defparam ram16s_inst_621.INIT_0 = 16'h0000;
defparam ram16s_inst_621.INIT_1 = 16'h8000;
defparam ram16s_inst_621.INIT_2 = 16'h07F0;
defparam ram16s_inst_621.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_622 (
    .DO(ram16s_inst_622_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2491),
    .CLK(clk)
);

defparam ram16s_inst_622.INIT_0 = 16'h0000;
defparam ram16s_inst_622.INIT_1 = 16'hFC3F;
defparam ram16s_inst_622.INIT_2 = 16'h0000;
defparam ram16s_inst_622.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_623 (
    .DO(ram16s_inst_623_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2495),
    .CLK(clk)
);

defparam ram16s_inst_623.INIT_0 = 16'h0000;
defparam ram16s_inst_623.INIT_1 = 16'h0001;
defparam ram16s_inst_623.INIT_2 = 16'h0000;
defparam ram16s_inst_623.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_624 (
    .DO(ram16s_inst_624_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2499),
    .CLK(clk)
);

defparam ram16s_inst_624.INIT_0 = 16'h0000;
defparam ram16s_inst_624.INIT_1 = 16'h0000;
defparam ram16s_inst_624.INIT_2 = 16'h0000;
defparam ram16s_inst_624.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_625 (
    .DO(ram16s_inst_625_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2503),
    .CLK(clk)
);

defparam ram16s_inst_625.INIT_0 = 16'h0000;
defparam ram16s_inst_625.INIT_1 = 16'h0000;
defparam ram16s_inst_625.INIT_2 = 16'hFE00;
defparam ram16s_inst_625.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_626 (
    .DO(ram16s_inst_626_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2507),
    .CLK(clk)
);

defparam ram16s_inst_626.INIT_0 = 16'h0000;
defparam ram16s_inst_626.INIT_1 = 16'h8000;
defparam ram16s_inst_626.INIT_2 = 16'h07F0;
defparam ram16s_inst_626.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_627 (
    .DO(ram16s_inst_627_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2511),
    .CLK(clk)
);

defparam ram16s_inst_627.INIT_0 = 16'h0000;
defparam ram16s_inst_627.INIT_1 = 16'hFC3F;
defparam ram16s_inst_627.INIT_2 = 16'h0000;
defparam ram16s_inst_627.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_628 (
    .DO(ram16s_inst_628_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2515),
    .CLK(clk)
);

defparam ram16s_inst_628.INIT_0 = 16'h0000;
defparam ram16s_inst_628.INIT_1 = 16'h0001;
defparam ram16s_inst_628.INIT_2 = 16'h0000;
defparam ram16s_inst_628.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_629 (
    .DO(ram16s_inst_629_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2519),
    .CLK(clk)
);

defparam ram16s_inst_629.INIT_0 = 16'h0000;
defparam ram16s_inst_629.INIT_1 = 16'h0000;
defparam ram16s_inst_629.INIT_2 = 16'h0000;
defparam ram16s_inst_629.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_630 (
    .DO(ram16s_inst_630_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2523),
    .CLK(clk)
);

defparam ram16s_inst_630.INIT_0 = 16'h0000;
defparam ram16s_inst_630.INIT_1 = 16'h0000;
defparam ram16s_inst_630.INIT_2 = 16'hFE00;
defparam ram16s_inst_630.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_631 (
    .DO(ram16s_inst_631_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2527),
    .CLK(clk)
);

defparam ram16s_inst_631.INIT_0 = 16'h0000;
defparam ram16s_inst_631.INIT_1 = 16'h8000;
defparam ram16s_inst_631.INIT_2 = 16'h07F0;
defparam ram16s_inst_631.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_632 (
    .DO(ram16s_inst_632_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2531),
    .CLK(clk)
);

defparam ram16s_inst_632.INIT_0 = 16'h0000;
defparam ram16s_inst_632.INIT_1 = 16'hFC3F;
defparam ram16s_inst_632.INIT_2 = 16'h0000;
defparam ram16s_inst_632.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_633 (
    .DO(ram16s_inst_633_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2535),
    .CLK(clk)
);

defparam ram16s_inst_633.INIT_0 = 16'h0000;
defparam ram16s_inst_633.INIT_1 = 16'h0001;
defparam ram16s_inst_633.INIT_2 = 16'h0000;
defparam ram16s_inst_633.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_634 (
    .DO(ram16s_inst_634_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2539),
    .CLK(clk)
);

defparam ram16s_inst_634.INIT_0 = 16'h0000;
defparam ram16s_inst_634.INIT_1 = 16'h0000;
defparam ram16s_inst_634.INIT_2 = 16'h0000;
defparam ram16s_inst_634.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_635 (
    .DO(ram16s_inst_635_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2543),
    .CLK(clk)
);

defparam ram16s_inst_635.INIT_0 = 16'h0000;
defparam ram16s_inst_635.INIT_1 = 16'h0000;
defparam ram16s_inst_635.INIT_2 = 16'hFE00;
defparam ram16s_inst_635.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_636 (
    .DO(ram16s_inst_636_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2547),
    .CLK(clk)
);

defparam ram16s_inst_636.INIT_0 = 16'h0000;
defparam ram16s_inst_636.INIT_1 = 16'h8000;
defparam ram16s_inst_636.INIT_2 = 16'h07F0;
defparam ram16s_inst_636.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_637 (
    .DO(ram16s_inst_637_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2551),
    .CLK(clk)
);

defparam ram16s_inst_637.INIT_0 = 16'h0000;
defparam ram16s_inst_637.INIT_1 = 16'hFC3F;
defparam ram16s_inst_637.INIT_2 = 16'h0000;
defparam ram16s_inst_637.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_638 (
    .DO(ram16s_inst_638_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2555),
    .CLK(clk)
);

defparam ram16s_inst_638.INIT_0 = 16'h0000;
defparam ram16s_inst_638.INIT_1 = 16'h0001;
defparam ram16s_inst_638.INIT_2 = 16'h0000;
defparam ram16s_inst_638.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_639 (
    .DO(ram16s_inst_639_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2559),
    .CLK(clk)
);

defparam ram16s_inst_639.INIT_0 = 16'h0000;
defparam ram16s_inst_639.INIT_1 = 16'h0000;
defparam ram16s_inst_639.INIT_2 = 16'h0000;
defparam ram16s_inst_639.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_640 (
    .DO(ram16s_inst_640_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2563),
    .CLK(clk)
);

defparam ram16s_inst_640.INIT_0 = 16'h0000;
defparam ram16s_inst_640.INIT_1 = 16'h0000;
defparam ram16s_inst_640.INIT_2 = 16'hFE00;
defparam ram16s_inst_640.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_641 (
    .DO(ram16s_inst_641_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2567),
    .CLK(clk)
);

defparam ram16s_inst_641.INIT_0 = 16'h0000;
defparam ram16s_inst_641.INIT_1 = 16'h8000;
defparam ram16s_inst_641.INIT_2 = 16'h07F0;
defparam ram16s_inst_641.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_642 (
    .DO(ram16s_inst_642_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2571),
    .CLK(clk)
);

defparam ram16s_inst_642.INIT_0 = 16'h0000;
defparam ram16s_inst_642.INIT_1 = 16'hFC3F;
defparam ram16s_inst_642.INIT_2 = 16'h0000;
defparam ram16s_inst_642.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_643 (
    .DO(ram16s_inst_643_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2575),
    .CLK(clk)
);

defparam ram16s_inst_643.INIT_0 = 16'h0000;
defparam ram16s_inst_643.INIT_1 = 16'h0001;
defparam ram16s_inst_643.INIT_2 = 16'h0000;
defparam ram16s_inst_643.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_644 (
    .DO(ram16s_inst_644_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2579),
    .CLK(clk)
);

defparam ram16s_inst_644.INIT_0 = 16'h0000;
defparam ram16s_inst_644.INIT_1 = 16'h0000;
defparam ram16s_inst_644.INIT_2 = 16'h0000;
defparam ram16s_inst_644.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_645 (
    .DO(ram16s_inst_645_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2583),
    .CLK(clk)
);

defparam ram16s_inst_645.INIT_0 = 16'h0000;
defparam ram16s_inst_645.INIT_1 = 16'h0000;
defparam ram16s_inst_645.INIT_2 = 16'h0000;
defparam ram16s_inst_645.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_646 (
    .DO(ram16s_inst_646_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2587),
    .CLK(clk)
);

defparam ram16s_inst_646.INIT_0 = 16'h0000;
defparam ram16s_inst_646.INIT_1 = 16'h0000;
defparam ram16s_inst_646.INIT_2 = 16'h0000;
defparam ram16s_inst_646.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_647 (
    .DO(ram16s_inst_647_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2591),
    .CLK(clk)
);

defparam ram16s_inst_647.INIT_0 = 16'h0000;
defparam ram16s_inst_647.INIT_1 = 16'h0000;
defparam ram16s_inst_647.INIT_2 = 16'h0000;
defparam ram16s_inst_647.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_648 (
    .DO(ram16s_inst_648_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2595),
    .CLK(clk)
);

defparam ram16s_inst_648.INIT_0 = 16'h0000;
defparam ram16s_inst_648.INIT_1 = 16'h0000;
defparam ram16s_inst_648.INIT_2 = 16'h0000;
defparam ram16s_inst_648.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_649 (
    .DO(ram16s_inst_649_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2599),
    .CLK(clk)
);

defparam ram16s_inst_649.INIT_0 = 16'h0000;
defparam ram16s_inst_649.INIT_1 = 16'h0000;
defparam ram16s_inst_649.INIT_2 = 16'h0000;
defparam ram16s_inst_649.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_650 (
    .DO(ram16s_inst_650_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2603),
    .CLK(clk)
);

defparam ram16s_inst_650.INIT_0 = 16'h0000;
defparam ram16s_inst_650.INIT_1 = 16'h0000;
defparam ram16s_inst_650.INIT_2 = 16'h0000;
defparam ram16s_inst_650.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_651 (
    .DO(ram16s_inst_651_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2607),
    .CLK(clk)
);

defparam ram16s_inst_651.INIT_0 = 16'h0000;
defparam ram16s_inst_651.INIT_1 = 16'h0000;
defparam ram16s_inst_651.INIT_2 = 16'h0000;
defparam ram16s_inst_651.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_652 (
    .DO(ram16s_inst_652_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2611),
    .CLK(clk)
);

defparam ram16s_inst_652.INIT_0 = 16'h0000;
defparam ram16s_inst_652.INIT_1 = 16'h0000;
defparam ram16s_inst_652.INIT_2 = 16'h0000;
defparam ram16s_inst_652.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_653 (
    .DO(ram16s_inst_653_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2615),
    .CLK(clk)
);

defparam ram16s_inst_653.INIT_0 = 16'h0000;
defparam ram16s_inst_653.INIT_1 = 16'h0000;
defparam ram16s_inst_653.INIT_2 = 16'h0000;
defparam ram16s_inst_653.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_654 (
    .DO(ram16s_inst_654_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2619),
    .CLK(clk)
);

defparam ram16s_inst_654.INIT_0 = 16'h0000;
defparam ram16s_inst_654.INIT_1 = 16'h0000;
defparam ram16s_inst_654.INIT_2 = 16'h0000;
defparam ram16s_inst_654.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_655 (
    .DO(ram16s_inst_655_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2623),
    .CLK(clk)
);

defparam ram16s_inst_655.INIT_0 = 16'h0000;
defparam ram16s_inst_655.INIT_1 = 16'h0000;
defparam ram16s_inst_655.INIT_2 = 16'h0000;
defparam ram16s_inst_655.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_656 (
    .DO(ram16s_inst_656_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2627),
    .CLK(clk)
);

defparam ram16s_inst_656.INIT_0 = 16'h0000;
defparam ram16s_inst_656.INIT_1 = 16'h0000;
defparam ram16s_inst_656.INIT_2 = 16'h0000;
defparam ram16s_inst_656.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_657 (
    .DO(ram16s_inst_657_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2631),
    .CLK(clk)
);

defparam ram16s_inst_657.INIT_0 = 16'h0000;
defparam ram16s_inst_657.INIT_1 = 16'h0000;
defparam ram16s_inst_657.INIT_2 = 16'h0000;
defparam ram16s_inst_657.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_658 (
    .DO(ram16s_inst_658_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2635),
    .CLK(clk)
);

defparam ram16s_inst_658.INIT_0 = 16'h0000;
defparam ram16s_inst_658.INIT_1 = 16'h0000;
defparam ram16s_inst_658.INIT_2 = 16'h0000;
defparam ram16s_inst_658.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_659 (
    .DO(ram16s_inst_659_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2639),
    .CLK(clk)
);

defparam ram16s_inst_659.INIT_0 = 16'h0000;
defparam ram16s_inst_659.INIT_1 = 16'h0000;
defparam ram16s_inst_659.INIT_2 = 16'h0000;
defparam ram16s_inst_659.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_660 (
    .DO(ram16s_inst_660_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2643),
    .CLK(clk)
);

defparam ram16s_inst_660.INIT_0 = 16'h0000;
defparam ram16s_inst_660.INIT_1 = 16'h0000;
defparam ram16s_inst_660.INIT_2 = 16'hFE00;
defparam ram16s_inst_660.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_661 (
    .DO(ram16s_inst_661_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2647),
    .CLK(clk)
);

defparam ram16s_inst_661.INIT_0 = 16'h0000;
defparam ram16s_inst_661.INIT_1 = 16'h8000;
defparam ram16s_inst_661.INIT_2 = 16'h07F0;
defparam ram16s_inst_661.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_662 (
    .DO(ram16s_inst_662_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2651),
    .CLK(clk)
);

defparam ram16s_inst_662.INIT_0 = 16'h0000;
defparam ram16s_inst_662.INIT_1 = 16'hFC3F;
defparam ram16s_inst_662.INIT_2 = 16'h0000;
defparam ram16s_inst_662.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_663 (
    .DO(ram16s_inst_663_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2655),
    .CLK(clk)
);

defparam ram16s_inst_663.INIT_0 = 16'h0000;
defparam ram16s_inst_663.INIT_1 = 16'h0001;
defparam ram16s_inst_663.INIT_2 = 16'h0000;
defparam ram16s_inst_663.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_664 (
    .DO(ram16s_inst_664_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2659),
    .CLK(clk)
);

defparam ram16s_inst_664.INIT_0 = 16'h0000;
defparam ram16s_inst_664.INIT_1 = 16'h0000;
defparam ram16s_inst_664.INIT_2 = 16'h0000;
defparam ram16s_inst_664.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_665 (
    .DO(ram16s_inst_665_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2663),
    .CLK(clk)
);

defparam ram16s_inst_665.INIT_0 = 16'h0000;
defparam ram16s_inst_665.INIT_1 = 16'h0000;
defparam ram16s_inst_665.INIT_2 = 16'hFE00;
defparam ram16s_inst_665.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_666 (
    .DO(ram16s_inst_666_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2667),
    .CLK(clk)
);

defparam ram16s_inst_666.INIT_0 = 16'h0000;
defparam ram16s_inst_666.INIT_1 = 16'h8000;
defparam ram16s_inst_666.INIT_2 = 16'h07F0;
defparam ram16s_inst_666.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_667 (
    .DO(ram16s_inst_667_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2671),
    .CLK(clk)
);

defparam ram16s_inst_667.INIT_0 = 16'h0000;
defparam ram16s_inst_667.INIT_1 = 16'hFC3F;
defparam ram16s_inst_667.INIT_2 = 16'h0000;
defparam ram16s_inst_667.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_668 (
    .DO(ram16s_inst_668_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2675),
    .CLK(clk)
);

defparam ram16s_inst_668.INIT_0 = 16'h0000;
defparam ram16s_inst_668.INIT_1 = 16'h0001;
defparam ram16s_inst_668.INIT_2 = 16'h0000;
defparam ram16s_inst_668.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_669 (
    .DO(ram16s_inst_669_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2679),
    .CLK(clk)
);

defparam ram16s_inst_669.INIT_0 = 16'h0000;
defparam ram16s_inst_669.INIT_1 = 16'h0000;
defparam ram16s_inst_669.INIT_2 = 16'h0000;
defparam ram16s_inst_669.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_670 (
    .DO(ram16s_inst_670_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2683),
    .CLK(clk)
);

defparam ram16s_inst_670.INIT_0 = 16'h0000;
defparam ram16s_inst_670.INIT_1 = 16'h0000;
defparam ram16s_inst_670.INIT_2 = 16'hFE00;
defparam ram16s_inst_670.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_671 (
    .DO(ram16s_inst_671_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2687),
    .CLK(clk)
);

defparam ram16s_inst_671.INIT_0 = 16'h0000;
defparam ram16s_inst_671.INIT_1 = 16'h8000;
defparam ram16s_inst_671.INIT_2 = 16'h07F0;
defparam ram16s_inst_671.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_672 (
    .DO(ram16s_inst_672_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2691),
    .CLK(clk)
);

defparam ram16s_inst_672.INIT_0 = 16'h0000;
defparam ram16s_inst_672.INIT_1 = 16'hFC3F;
defparam ram16s_inst_672.INIT_2 = 16'h0000;
defparam ram16s_inst_672.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_673 (
    .DO(ram16s_inst_673_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2695),
    .CLK(clk)
);

defparam ram16s_inst_673.INIT_0 = 16'h0000;
defparam ram16s_inst_673.INIT_1 = 16'h0001;
defparam ram16s_inst_673.INIT_2 = 16'h0000;
defparam ram16s_inst_673.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_674 (
    .DO(ram16s_inst_674_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2699),
    .CLK(clk)
);

defparam ram16s_inst_674.INIT_0 = 16'h0000;
defparam ram16s_inst_674.INIT_1 = 16'h0000;
defparam ram16s_inst_674.INIT_2 = 16'h0000;
defparam ram16s_inst_674.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_675 (
    .DO(ram16s_inst_675_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2703),
    .CLK(clk)
);

defparam ram16s_inst_675.INIT_0 = 16'h0000;
defparam ram16s_inst_675.INIT_1 = 16'h0000;
defparam ram16s_inst_675.INIT_2 = 16'hFE00;
defparam ram16s_inst_675.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_676 (
    .DO(ram16s_inst_676_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2707),
    .CLK(clk)
);

defparam ram16s_inst_676.INIT_0 = 16'h0000;
defparam ram16s_inst_676.INIT_1 = 16'h8000;
defparam ram16s_inst_676.INIT_2 = 16'h07F0;
defparam ram16s_inst_676.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_677 (
    .DO(ram16s_inst_677_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2711),
    .CLK(clk)
);

defparam ram16s_inst_677.INIT_0 = 16'h0000;
defparam ram16s_inst_677.INIT_1 = 16'hFC3F;
defparam ram16s_inst_677.INIT_2 = 16'h0000;
defparam ram16s_inst_677.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_678 (
    .DO(ram16s_inst_678_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2715),
    .CLK(clk)
);

defparam ram16s_inst_678.INIT_0 = 16'h0000;
defparam ram16s_inst_678.INIT_1 = 16'h0001;
defparam ram16s_inst_678.INIT_2 = 16'h0000;
defparam ram16s_inst_678.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_679 (
    .DO(ram16s_inst_679_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2719),
    .CLK(clk)
);

defparam ram16s_inst_679.INIT_0 = 16'h0000;
defparam ram16s_inst_679.INIT_1 = 16'h0000;
defparam ram16s_inst_679.INIT_2 = 16'h0000;
defparam ram16s_inst_679.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_680 (
    .DO(ram16s_inst_680_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2723),
    .CLK(clk)
);

defparam ram16s_inst_680.INIT_0 = 16'h0000;
defparam ram16s_inst_680.INIT_1 = 16'h0000;
defparam ram16s_inst_680.INIT_2 = 16'hFE00;
defparam ram16s_inst_680.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_681 (
    .DO(ram16s_inst_681_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2727),
    .CLK(clk)
);

defparam ram16s_inst_681.INIT_0 = 16'h0000;
defparam ram16s_inst_681.INIT_1 = 16'h8000;
defparam ram16s_inst_681.INIT_2 = 16'h07F0;
defparam ram16s_inst_681.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_682 (
    .DO(ram16s_inst_682_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2731),
    .CLK(clk)
);

defparam ram16s_inst_682.INIT_0 = 16'h0000;
defparam ram16s_inst_682.INIT_1 = 16'hFC3F;
defparam ram16s_inst_682.INIT_2 = 16'h0000;
defparam ram16s_inst_682.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_683 (
    .DO(ram16s_inst_683_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2735),
    .CLK(clk)
);

defparam ram16s_inst_683.INIT_0 = 16'h0000;
defparam ram16s_inst_683.INIT_1 = 16'h0001;
defparam ram16s_inst_683.INIT_2 = 16'h0000;
defparam ram16s_inst_683.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_684 (
    .DO(ram16s_inst_684_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2739),
    .CLK(clk)
);

defparam ram16s_inst_684.INIT_0 = 16'h0000;
defparam ram16s_inst_684.INIT_1 = 16'h0000;
defparam ram16s_inst_684.INIT_2 = 16'h0000;
defparam ram16s_inst_684.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_685 (
    .DO(ram16s_inst_685_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2743),
    .CLK(clk)
);

defparam ram16s_inst_685.INIT_0 = 16'h0000;
defparam ram16s_inst_685.INIT_1 = 16'h0000;
defparam ram16s_inst_685.INIT_2 = 16'hFE00;
defparam ram16s_inst_685.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_686 (
    .DO(ram16s_inst_686_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2747),
    .CLK(clk)
);

defparam ram16s_inst_686.INIT_0 = 16'h0000;
defparam ram16s_inst_686.INIT_1 = 16'h8000;
defparam ram16s_inst_686.INIT_2 = 16'h07F0;
defparam ram16s_inst_686.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_687 (
    .DO(ram16s_inst_687_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2751),
    .CLK(clk)
);

defparam ram16s_inst_687.INIT_0 = 16'h0000;
defparam ram16s_inst_687.INIT_1 = 16'hFC3F;
defparam ram16s_inst_687.INIT_2 = 16'h0000;
defparam ram16s_inst_687.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_688 (
    .DO(ram16s_inst_688_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2755),
    .CLK(clk)
);

defparam ram16s_inst_688.INIT_0 = 16'h0000;
defparam ram16s_inst_688.INIT_1 = 16'h0001;
defparam ram16s_inst_688.INIT_2 = 16'h0000;
defparam ram16s_inst_688.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_689 (
    .DO(ram16s_inst_689_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2759),
    .CLK(clk)
);

defparam ram16s_inst_689.INIT_0 = 16'h0000;
defparam ram16s_inst_689.INIT_1 = 16'h0000;
defparam ram16s_inst_689.INIT_2 = 16'h0000;
defparam ram16s_inst_689.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_690 (
    .DO(ram16s_inst_690_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2763),
    .CLK(clk)
);

defparam ram16s_inst_690.INIT_0 = 16'h0000;
defparam ram16s_inst_690.INIT_1 = 16'h0000;
defparam ram16s_inst_690.INIT_2 = 16'h0000;
defparam ram16s_inst_690.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_691 (
    .DO(ram16s_inst_691_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2767),
    .CLK(clk)
);

defparam ram16s_inst_691.INIT_0 = 16'h0000;
defparam ram16s_inst_691.INIT_1 = 16'h0000;
defparam ram16s_inst_691.INIT_2 = 16'h0000;
defparam ram16s_inst_691.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_692 (
    .DO(ram16s_inst_692_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2771),
    .CLK(clk)
);

defparam ram16s_inst_692.INIT_0 = 16'h0000;
defparam ram16s_inst_692.INIT_1 = 16'h0000;
defparam ram16s_inst_692.INIT_2 = 16'h0000;
defparam ram16s_inst_692.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_693 (
    .DO(ram16s_inst_693_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2775),
    .CLK(clk)
);

defparam ram16s_inst_693.INIT_0 = 16'h0000;
defparam ram16s_inst_693.INIT_1 = 16'h0000;
defparam ram16s_inst_693.INIT_2 = 16'h0000;
defparam ram16s_inst_693.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_694 (
    .DO(ram16s_inst_694_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2779),
    .CLK(clk)
);

defparam ram16s_inst_694.INIT_0 = 16'h0000;
defparam ram16s_inst_694.INIT_1 = 16'h0000;
defparam ram16s_inst_694.INIT_2 = 16'h0000;
defparam ram16s_inst_694.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_695 (
    .DO(ram16s_inst_695_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2783),
    .CLK(clk)
);

defparam ram16s_inst_695.INIT_0 = 16'h0000;
defparam ram16s_inst_695.INIT_1 = 16'h0000;
defparam ram16s_inst_695.INIT_2 = 16'h0000;
defparam ram16s_inst_695.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_696 (
    .DO(ram16s_inst_696_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2787),
    .CLK(clk)
);

defparam ram16s_inst_696.INIT_0 = 16'h0000;
defparam ram16s_inst_696.INIT_1 = 16'h0000;
defparam ram16s_inst_696.INIT_2 = 16'h0000;
defparam ram16s_inst_696.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_697 (
    .DO(ram16s_inst_697_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2791),
    .CLK(clk)
);

defparam ram16s_inst_697.INIT_0 = 16'h0000;
defparam ram16s_inst_697.INIT_1 = 16'h0000;
defparam ram16s_inst_697.INIT_2 = 16'h0000;
defparam ram16s_inst_697.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_698 (
    .DO(ram16s_inst_698_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2795),
    .CLK(clk)
);

defparam ram16s_inst_698.INIT_0 = 16'h0000;
defparam ram16s_inst_698.INIT_1 = 16'h0000;
defparam ram16s_inst_698.INIT_2 = 16'h0000;
defparam ram16s_inst_698.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_699 (
    .DO(ram16s_inst_699_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2799),
    .CLK(clk)
);

defparam ram16s_inst_699.INIT_0 = 16'h0000;
defparam ram16s_inst_699.INIT_1 = 16'h0000;
defparam ram16s_inst_699.INIT_2 = 16'h0000;
defparam ram16s_inst_699.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_700 (
    .DO(ram16s_inst_700_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2803),
    .CLK(clk)
);

defparam ram16s_inst_700.INIT_0 = 16'h0000;
defparam ram16s_inst_700.INIT_1 = 16'h0000;
defparam ram16s_inst_700.INIT_2 = 16'h0000;
defparam ram16s_inst_700.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_701 (
    .DO(ram16s_inst_701_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2807),
    .CLK(clk)
);

defparam ram16s_inst_701.INIT_0 = 16'h0000;
defparam ram16s_inst_701.INIT_1 = 16'h0000;
defparam ram16s_inst_701.INIT_2 = 16'h0000;
defparam ram16s_inst_701.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_702 (
    .DO(ram16s_inst_702_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2811),
    .CLK(clk)
);

defparam ram16s_inst_702.INIT_0 = 16'h0000;
defparam ram16s_inst_702.INIT_1 = 16'h0000;
defparam ram16s_inst_702.INIT_2 = 16'h0000;
defparam ram16s_inst_702.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_703 (
    .DO(ram16s_inst_703_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2815),
    .CLK(clk)
);

defparam ram16s_inst_703.INIT_0 = 16'h0000;
defparam ram16s_inst_703.INIT_1 = 16'h0000;
defparam ram16s_inst_703.INIT_2 = 16'h0000;
defparam ram16s_inst_703.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_704 (
    .DO(ram16s_inst_704_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2819),
    .CLK(clk)
);

defparam ram16s_inst_704.INIT_0 = 16'h0000;
defparam ram16s_inst_704.INIT_1 = 16'h0000;
defparam ram16s_inst_704.INIT_2 = 16'h0000;
defparam ram16s_inst_704.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_705 (
    .DO(ram16s_inst_705_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2823),
    .CLK(clk)
);

defparam ram16s_inst_705.INIT_0 = 16'h0000;
defparam ram16s_inst_705.INIT_1 = 16'h0000;
defparam ram16s_inst_705.INIT_2 = 16'h0000;
defparam ram16s_inst_705.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_706 (
    .DO(ram16s_inst_706_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2827),
    .CLK(clk)
);

defparam ram16s_inst_706.INIT_0 = 16'h0000;
defparam ram16s_inst_706.INIT_1 = 16'h0000;
defparam ram16s_inst_706.INIT_2 = 16'h0000;
defparam ram16s_inst_706.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_707 (
    .DO(ram16s_inst_707_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2831),
    .CLK(clk)
);

defparam ram16s_inst_707.INIT_0 = 16'h0000;
defparam ram16s_inst_707.INIT_1 = 16'h0000;
defparam ram16s_inst_707.INIT_2 = 16'h0000;
defparam ram16s_inst_707.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_708 (
    .DO(ram16s_inst_708_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2835),
    .CLK(clk)
);

defparam ram16s_inst_708.INIT_0 = 16'h0000;
defparam ram16s_inst_708.INIT_1 = 16'h0000;
defparam ram16s_inst_708.INIT_2 = 16'h0000;
defparam ram16s_inst_708.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_709 (
    .DO(ram16s_inst_709_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2839),
    .CLK(clk)
);

defparam ram16s_inst_709.INIT_0 = 16'h0000;
defparam ram16s_inst_709.INIT_1 = 16'h0000;
defparam ram16s_inst_709.INIT_2 = 16'h0000;
defparam ram16s_inst_709.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_710 (
    .DO(ram16s_inst_710_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2843),
    .CLK(clk)
);

defparam ram16s_inst_710.INIT_0 = 16'h0000;
defparam ram16s_inst_710.INIT_1 = 16'h0000;
defparam ram16s_inst_710.INIT_2 = 16'h0000;
defparam ram16s_inst_710.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_711 (
    .DO(ram16s_inst_711_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2847),
    .CLK(clk)
);

defparam ram16s_inst_711.INIT_0 = 16'h0000;
defparam ram16s_inst_711.INIT_1 = 16'h0000;
defparam ram16s_inst_711.INIT_2 = 16'h0000;
defparam ram16s_inst_711.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_712 (
    .DO(ram16s_inst_712_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2851),
    .CLK(clk)
);

defparam ram16s_inst_712.INIT_0 = 16'h0000;
defparam ram16s_inst_712.INIT_1 = 16'h0000;
defparam ram16s_inst_712.INIT_2 = 16'h0000;
defparam ram16s_inst_712.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_713 (
    .DO(ram16s_inst_713_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2855),
    .CLK(clk)
);

defparam ram16s_inst_713.INIT_0 = 16'h0000;
defparam ram16s_inst_713.INIT_1 = 16'h0000;
defparam ram16s_inst_713.INIT_2 = 16'h0000;
defparam ram16s_inst_713.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_714 (
    .DO(ram16s_inst_714_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2859),
    .CLK(clk)
);

defparam ram16s_inst_714.INIT_0 = 16'h0000;
defparam ram16s_inst_714.INIT_1 = 16'h0000;
defparam ram16s_inst_714.INIT_2 = 16'h0000;
defparam ram16s_inst_714.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_715 (
    .DO(ram16s_inst_715_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2863),
    .CLK(clk)
);

defparam ram16s_inst_715.INIT_0 = 16'h0000;
defparam ram16s_inst_715.INIT_1 = 16'h0000;
defparam ram16s_inst_715.INIT_2 = 16'h0000;
defparam ram16s_inst_715.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_716 (
    .DO(ram16s_inst_716_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2867),
    .CLK(clk)
);

defparam ram16s_inst_716.INIT_0 = 16'h0000;
defparam ram16s_inst_716.INIT_1 = 16'h0000;
defparam ram16s_inst_716.INIT_2 = 16'h0000;
defparam ram16s_inst_716.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_717 (
    .DO(ram16s_inst_717_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2871),
    .CLK(clk)
);

defparam ram16s_inst_717.INIT_0 = 16'h0000;
defparam ram16s_inst_717.INIT_1 = 16'h0000;
defparam ram16s_inst_717.INIT_2 = 16'h0000;
defparam ram16s_inst_717.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_718 (
    .DO(ram16s_inst_718_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2875),
    .CLK(clk)
);

defparam ram16s_inst_718.INIT_0 = 16'h0000;
defparam ram16s_inst_718.INIT_1 = 16'h0000;
defparam ram16s_inst_718.INIT_2 = 16'h0000;
defparam ram16s_inst_718.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_719 (
    .DO(ram16s_inst_719_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2879),
    .CLK(clk)
);

defparam ram16s_inst_719.INIT_0 = 16'h0000;
defparam ram16s_inst_719.INIT_1 = 16'h0000;
defparam ram16s_inst_719.INIT_2 = 16'h0000;
defparam ram16s_inst_719.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_720 (
    .DO(ram16s_inst_720_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2883),
    .CLK(clk)
);

defparam ram16s_inst_720.INIT_0 = 16'h0000;
defparam ram16s_inst_720.INIT_1 = 16'h0000;
defparam ram16s_inst_720.INIT_2 = 16'h0000;
defparam ram16s_inst_720.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_721 (
    .DO(ram16s_inst_721_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2887),
    .CLK(clk)
);

defparam ram16s_inst_721.INIT_0 = 16'h0000;
defparam ram16s_inst_721.INIT_1 = 16'h0000;
defparam ram16s_inst_721.INIT_2 = 16'h0000;
defparam ram16s_inst_721.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_722 (
    .DO(ram16s_inst_722_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2891),
    .CLK(clk)
);

defparam ram16s_inst_722.INIT_0 = 16'h0000;
defparam ram16s_inst_722.INIT_1 = 16'h0000;
defparam ram16s_inst_722.INIT_2 = 16'h0000;
defparam ram16s_inst_722.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_723 (
    .DO(ram16s_inst_723_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2895),
    .CLK(clk)
);

defparam ram16s_inst_723.INIT_0 = 16'h0000;
defparam ram16s_inst_723.INIT_1 = 16'h0000;
defparam ram16s_inst_723.INIT_2 = 16'h0000;
defparam ram16s_inst_723.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_724 (
    .DO(ram16s_inst_724_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2899),
    .CLK(clk)
);

defparam ram16s_inst_724.INIT_0 = 16'h0000;
defparam ram16s_inst_724.INIT_1 = 16'h0000;
defparam ram16s_inst_724.INIT_2 = 16'h0000;
defparam ram16s_inst_724.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_725 (
    .DO(ram16s_inst_725_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2903),
    .CLK(clk)
);

defparam ram16s_inst_725.INIT_0 = 16'h0000;
defparam ram16s_inst_725.INIT_1 = 16'h0000;
defparam ram16s_inst_725.INIT_2 = 16'h0000;
defparam ram16s_inst_725.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_726 (
    .DO(ram16s_inst_726_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2907),
    .CLK(clk)
);

defparam ram16s_inst_726.INIT_0 = 16'h0000;
defparam ram16s_inst_726.INIT_1 = 16'h0000;
defparam ram16s_inst_726.INIT_2 = 16'h0000;
defparam ram16s_inst_726.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_727 (
    .DO(ram16s_inst_727_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2911),
    .CLK(clk)
);

defparam ram16s_inst_727.INIT_0 = 16'h0000;
defparam ram16s_inst_727.INIT_1 = 16'h0000;
defparam ram16s_inst_727.INIT_2 = 16'h0000;
defparam ram16s_inst_727.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_728 (
    .DO(ram16s_inst_728_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2915),
    .CLK(clk)
);

defparam ram16s_inst_728.INIT_0 = 16'h0000;
defparam ram16s_inst_728.INIT_1 = 16'h0000;
defparam ram16s_inst_728.INIT_2 = 16'h0000;
defparam ram16s_inst_728.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_729 (
    .DO(ram16s_inst_729_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2919),
    .CLK(clk)
);

defparam ram16s_inst_729.INIT_0 = 16'h0000;
defparam ram16s_inst_729.INIT_1 = 16'h0000;
defparam ram16s_inst_729.INIT_2 = 16'h0000;
defparam ram16s_inst_729.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_730 (
    .DO(ram16s_inst_730_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2923),
    .CLK(clk)
);

defparam ram16s_inst_730.INIT_0 = 16'h0000;
defparam ram16s_inst_730.INIT_1 = 16'h0000;
defparam ram16s_inst_730.INIT_2 = 16'h0000;
defparam ram16s_inst_730.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_731 (
    .DO(ram16s_inst_731_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2927),
    .CLK(clk)
);

defparam ram16s_inst_731.INIT_0 = 16'h0000;
defparam ram16s_inst_731.INIT_1 = 16'h0000;
defparam ram16s_inst_731.INIT_2 = 16'h0000;
defparam ram16s_inst_731.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_732 (
    .DO(ram16s_inst_732_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2931),
    .CLK(clk)
);

defparam ram16s_inst_732.INIT_0 = 16'h0000;
defparam ram16s_inst_732.INIT_1 = 16'h0000;
defparam ram16s_inst_732.INIT_2 = 16'h0000;
defparam ram16s_inst_732.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_733 (
    .DO(ram16s_inst_733_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2935),
    .CLK(clk)
);

defparam ram16s_inst_733.INIT_0 = 16'h0000;
defparam ram16s_inst_733.INIT_1 = 16'h0000;
defparam ram16s_inst_733.INIT_2 = 16'h0000;
defparam ram16s_inst_733.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_734 (
    .DO(ram16s_inst_734_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2939),
    .CLK(clk)
);

defparam ram16s_inst_734.INIT_0 = 16'h0000;
defparam ram16s_inst_734.INIT_1 = 16'h0000;
defparam ram16s_inst_734.INIT_2 = 16'h0000;
defparam ram16s_inst_734.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_735 (
    .DO(ram16s_inst_735_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2943),
    .CLK(clk)
);

defparam ram16s_inst_735.INIT_0 = 16'h0000;
defparam ram16s_inst_735.INIT_1 = 16'h0000;
defparam ram16s_inst_735.INIT_2 = 16'h0000;
defparam ram16s_inst_735.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_736 (
    .DO(ram16s_inst_736_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2947),
    .CLK(clk)
);

defparam ram16s_inst_736.INIT_0 = 16'h0000;
defparam ram16s_inst_736.INIT_1 = 16'h0000;
defparam ram16s_inst_736.INIT_2 = 16'h0000;
defparam ram16s_inst_736.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_737 (
    .DO(ram16s_inst_737_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2951),
    .CLK(clk)
);

defparam ram16s_inst_737.INIT_0 = 16'h0000;
defparam ram16s_inst_737.INIT_1 = 16'h0000;
defparam ram16s_inst_737.INIT_2 = 16'h0000;
defparam ram16s_inst_737.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_738 (
    .DO(ram16s_inst_738_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2955),
    .CLK(clk)
);

defparam ram16s_inst_738.INIT_0 = 16'h0000;
defparam ram16s_inst_738.INIT_1 = 16'h0000;
defparam ram16s_inst_738.INIT_2 = 16'h0000;
defparam ram16s_inst_738.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_739 (
    .DO(ram16s_inst_739_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2959),
    .CLK(clk)
);

defparam ram16s_inst_739.INIT_0 = 16'h0000;
defparam ram16s_inst_739.INIT_1 = 16'h0000;
defparam ram16s_inst_739.INIT_2 = 16'h0000;
defparam ram16s_inst_739.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_740 (
    .DO(ram16s_inst_740_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2963),
    .CLK(clk)
);

defparam ram16s_inst_740.INIT_0 = 16'h0000;
defparam ram16s_inst_740.INIT_1 = 16'h0000;
defparam ram16s_inst_740.INIT_2 = 16'h0000;
defparam ram16s_inst_740.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_741 (
    .DO(ram16s_inst_741_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2967),
    .CLK(clk)
);

defparam ram16s_inst_741.INIT_0 = 16'h0000;
defparam ram16s_inst_741.INIT_1 = 16'h0000;
defparam ram16s_inst_741.INIT_2 = 16'h0000;
defparam ram16s_inst_741.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_742 (
    .DO(ram16s_inst_742_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2971),
    .CLK(clk)
);

defparam ram16s_inst_742.INIT_0 = 16'h0000;
defparam ram16s_inst_742.INIT_1 = 16'h0000;
defparam ram16s_inst_742.INIT_2 = 16'h0000;
defparam ram16s_inst_742.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_743 (
    .DO(ram16s_inst_743_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2975),
    .CLK(clk)
);

defparam ram16s_inst_743.INIT_0 = 16'h0000;
defparam ram16s_inst_743.INIT_1 = 16'h0000;
defparam ram16s_inst_743.INIT_2 = 16'h0000;
defparam ram16s_inst_743.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_744 (
    .DO(ram16s_inst_744_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2979),
    .CLK(clk)
);

defparam ram16s_inst_744.INIT_0 = 16'h0000;
defparam ram16s_inst_744.INIT_1 = 16'h0000;
defparam ram16s_inst_744.INIT_2 = 16'h0000;
defparam ram16s_inst_744.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_745 (
    .DO(ram16s_inst_745_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2983),
    .CLK(clk)
);

defparam ram16s_inst_745.INIT_0 = 16'h0000;
defparam ram16s_inst_745.INIT_1 = 16'h0000;
defparam ram16s_inst_745.INIT_2 = 16'h0000;
defparam ram16s_inst_745.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_746 (
    .DO(ram16s_inst_746_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2987),
    .CLK(clk)
);

defparam ram16s_inst_746.INIT_0 = 16'h0000;
defparam ram16s_inst_746.INIT_1 = 16'h0000;
defparam ram16s_inst_746.INIT_2 = 16'h0000;
defparam ram16s_inst_746.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_747 (
    .DO(ram16s_inst_747_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2991),
    .CLK(clk)
);

defparam ram16s_inst_747.INIT_0 = 16'h0000;
defparam ram16s_inst_747.INIT_1 = 16'h0000;
defparam ram16s_inst_747.INIT_2 = 16'h0000;
defparam ram16s_inst_747.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_748 (
    .DO(ram16s_inst_748_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2995),
    .CLK(clk)
);

defparam ram16s_inst_748.INIT_0 = 16'h0000;
defparam ram16s_inst_748.INIT_1 = 16'h0000;
defparam ram16s_inst_748.INIT_2 = 16'h0000;
defparam ram16s_inst_748.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_749 (
    .DO(ram16s_inst_749_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_2999),
    .CLK(clk)
);

defparam ram16s_inst_749.INIT_0 = 16'h0000;
defparam ram16s_inst_749.INIT_1 = 16'h0000;
defparam ram16s_inst_749.INIT_2 = 16'h0000;
defparam ram16s_inst_749.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_750 (
    .DO(ram16s_inst_750_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3003),
    .CLK(clk)
);

defparam ram16s_inst_750.INIT_0 = 16'h0000;
defparam ram16s_inst_750.INIT_1 = 16'h0000;
defparam ram16s_inst_750.INIT_2 = 16'h0000;
defparam ram16s_inst_750.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_751 (
    .DO(ram16s_inst_751_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3007),
    .CLK(clk)
);

defparam ram16s_inst_751.INIT_0 = 16'h0000;
defparam ram16s_inst_751.INIT_1 = 16'h0000;
defparam ram16s_inst_751.INIT_2 = 16'h0000;
defparam ram16s_inst_751.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_752 (
    .DO(ram16s_inst_752_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3011),
    .CLK(clk)
);

defparam ram16s_inst_752.INIT_0 = 16'h0000;
defparam ram16s_inst_752.INIT_1 = 16'h0000;
defparam ram16s_inst_752.INIT_2 = 16'h0000;
defparam ram16s_inst_752.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_753 (
    .DO(ram16s_inst_753_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3015),
    .CLK(clk)
);

defparam ram16s_inst_753.INIT_0 = 16'h0000;
defparam ram16s_inst_753.INIT_1 = 16'h0000;
defparam ram16s_inst_753.INIT_2 = 16'h0000;
defparam ram16s_inst_753.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_754 (
    .DO(ram16s_inst_754_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3019),
    .CLK(clk)
);

defparam ram16s_inst_754.INIT_0 = 16'h0000;
defparam ram16s_inst_754.INIT_1 = 16'h0000;
defparam ram16s_inst_754.INIT_2 = 16'h0000;
defparam ram16s_inst_754.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_755 (
    .DO(ram16s_inst_755_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3023),
    .CLK(clk)
);

defparam ram16s_inst_755.INIT_0 = 16'h0000;
defparam ram16s_inst_755.INIT_1 = 16'h0000;
defparam ram16s_inst_755.INIT_2 = 16'h0000;
defparam ram16s_inst_755.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_756 (
    .DO(ram16s_inst_756_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3027),
    .CLK(clk)
);

defparam ram16s_inst_756.INIT_0 = 16'h0000;
defparam ram16s_inst_756.INIT_1 = 16'h0000;
defparam ram16s_inst_756.INIT_2 = 16'h0000;
defparam ram16s_inst_756.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_757 (
    .DO(ram16s_inst_757_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3031),
    .CLK(clk)
);

defparam ram16s_inst_757.INIT_0 = 16'h0000;
defparam ram16s_inst_757.INIT_1 = 16'h0000;
defparam ram16s_inst_757.INIT_2 = 16'h0000;
defparam ram16s_inst_757.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_758 (
    .DO(ram16s_inst_758_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3035),
    .CLK(clk)
);

defparam ram16s_inst_758.INIT_0 = 16'h0000;
defparam ram16s_inst_758.INIT_1 = 16'h0000;
defparam ram16s_inst_758.INIT_2 = 16'h0000;
defparam ram16s_inst_758.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_759 (
    .DO(ram16s_inst_759_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3039),
    .CLK(clk)
);

defparam ram16s_inst_759.INIT_0 = 16'h0000;
defparam ram16s_inst_759.INIT_1 = 16'h0000;
defparam ram16s_inst_759.INIT_2 = 16'h0000;
defparam ram16s_inst_759.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_760 (
    .DO(ram16s_inst_760_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3043),
    .CLK(clk)
);

defparam ram16s_inst_760.INIT_0 = 16'h0000;
defparam ram16s_inst_760.INIT_1 = 16'h0000;
defparam ram16s_inst_760.INIT_2 = 16'h0000;
defparam ram16s_inst_760.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_761 (
    .DO(ram16s_inst_761_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3047),
    .CLK(clk)
);

defparam ram16s_inst_761.INIT_0 = 16'h0000;
defparam ram16s_inst_761.INIT_1 = 16'h0000;
defparam ram16s_inst_761.INIT_2 = 16'h0000;
defparam ram16s_inst_761.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_762 (
    .DO(ram16s_inst_762_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3051),
    .CLK(clk)
);

defparam ram16s_inst_762.INIT_0 = 16'h0000;
defparam ram16s_inst_762.INIT_1 = 16'h0000;
defparam ram16s_inst_762.INIT_2 = 16'h0000;
defparam ram16s_inst_762.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_763 (
    .DO(ram16s_inst_763_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3055),
    .CLK(clk)
);

defparam ram16s_inst_763.INIT_0 = 16'h0000;
defparam ram16s_inst_763.INIT_1 = 16'h0000;
defparam ram16s_inst_763.INIT_2 = 16'h0000;
defparam ram16s_inst_763.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_764 (
    .DO(ram16s_inst_764_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3059),
    .CLK(clk)
);

defparam ram16s_inst_764.INIT_0 = 16'h0000;
defparam ram16s_inst_764.INIT_1 = 16'h0000;
defparam ram16s_inst_764.INIT_2 = 16'h0000;
defparam ram16s_inst_764.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_765 (
    .DO(ram16s_inst_765_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3063),
    .CLK(clk)
);

defparam ram16s_inst_765.INIT_0 = 16'h0000;
defparam ram16s_inst_765.INIT_1 = 16'h0000;
defparam ram16s_inst_765.INIT_2 = 16'h0000;
defparam ram16s_inst_765.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_766 (
    .DO(ram16s_inst_766_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3067),
    .CLK(clk)
);

defparam ram16s_inst_766.INIT_0 = 16'h0000;
defparam ram16s_inst_766.INIT_1 = 16'h0000;
defparam ram16s_inst_766.INIT_2 = 16'h0000;
defparam ram16s_inst_766.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_767 (
    .DO(ram16s_inst_767_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3071),
    .CLK(clk)
);

defparam ram16s_inst_767.INIT_0 = 16'h0000;
defparam ram16s_inst_767.INIT_1 = 16'h0000;
defparam ram16s_inst_767.INIT_2 = 16'h0000;
defparam ram16s_inst_767.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_768 (
    .DO(ram16s_inst_768_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3075),
    .CLK(clk)
);

defparam ram16s_inst_768.INIT_0 = 16'h0000;
defparam ram16s_inst_768.INIT_1 = 16'h0000;
defparam ram16s_inst_768.INIT_2 = 16'h0000;
defparam ram16s_inst_768.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_769 (
    .DO(ram16s_inst_769_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3079),
    .CLK(clk)
);

defparam ram16s_inst_769.INIT_0 = 16'h0000;
defparam ram16s_inst_769.INIT_1 = 16'h0000;
defparam ram16s_inst_769.INIT_2 = 16'h0000;
defparam ram16s_inst_769.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_770 (
    .DO(ram16s_inst_770_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3083),
    .CLK(clk)
);

defparam ram16s_inst_770.INIT_0 = 16'h0000;
defparam ram16s_inst_770.INIT_1 = 16'h0000;
defparam ram16s_inst_770.INIT_2 = 16'h0000;
defparam ram16s_inst_770.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_771 (
    .DO(ram16s_inst_771_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3087),
    .CLK(clk)
);

defparam ram16s_inst_771.INIT_0 = 16'h0000;
defparam ram16s_inst_771.INIT_1 = 16'h0000;
defparam ram16s_inst_771.INIT_2 = 16'h0000;
defparam ram16s_inst_771.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_772 (
    .DO(ram16s_inst_772_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3091),
    .CLK(clk)
);

defparam ram16s_inst_772.INIT_0 = 16'h0000;
defparam ram16s_inst_772.INIT_1 = 16'h0000;
defparam ram16s_inst_772.INIT_2 = 16'h0000;
defparam ram16s_inst_772.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_773 (
    .DO(ram16s_inst_773_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3095),
    .CLK(clk)
);

defparam ram16s_inst_773.INIT_0 = 16'h0000;
defparam ram16s_inst_773.INIT_1 = 16'h0000;
defparam ram16s_inst_773.INIT_2 = 16'h0000;
defparam ram16s_inst_773.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_774 (
    .DO(ram16s_inst_774_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3099),
    .CLK(clk)
);

defparam ram16s_inst_774.INIT_0 = 16'h0000;
defparam ram16s_inst_774.INIT_1 = 16'h0000;
defparam ram16s_inst_774.INIT_2 = 16'h0000;
defparam ram16s_inst_774.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_775 (
    .DO(ram16s_inst_775_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3103),
    .CLK(clk)
);

defparam ram16s_inst_775.INIT_0 = 16'h0000;
defparam ram16s_inst_775.INIT_1 = 16'h0000;
defparam ram16s_inst_775.INIT_2 = 16'h0000;
defparam ram16s_inst_775.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_776 (
    .DO(ram16s_inst_776_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3107),
    .CLK(clk)
);

defparam ram16s_inst_776.INIT_0 = 16'h0000;
defparam ram16s_inst_776.INIT_1 = 16'h0000;
defparam ram16s_inst_776.INIT_2 = 16'h0000;
defparam ram16s_inst_776.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_777 (
    .DO(ram16s_inst_777_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3111),
    .CLK(clk)
);

defparam ram16s_inst_777.INIT_0 = 16'h0000;
defparam ram16s_inst_777.INIT_1 = 16'h0000;
defparam ram16s_inst_777.INIT_2 = 16'h0000;
defparam ram16s_inst_777.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_778 (
    .DO(ram16s_inst_778_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3115),
    .CLK(clk)
);

defparam ram16s_inst_778.INIT_0 = 16'h0000;
defparam ram16s_inst_778.INIT_1 = 16'h0000;
defparam ram16s_inst_778.INIT_2 = 16'h0000;
defparam ram16s_inst_778.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_779 (
    .DO(ram16s_inst_779_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3119),
    .CLK(clk)
);

defparam ram16s_inst_779.INIT_0 = 16'h0000;
defparam ram16s_inst_779.INIT_1 = 16'h0000;
defparam ram16s_inst_779.INIT_2 = 16'h0000;
defparam ram16s_inst_779.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_780 (
    .DO(ram16s_inst_780_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3123),
    .CLK(clk)
);

defparam ram16s_inst_780.INIT_0 = 16'h0000;
defparam ram16s_inst_780.INIT_1 = 16'h0000;
defparam ram16s_inst_780.INIT_2 = 16'h0000;
defparam ram16s_inst_780.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_781 (
    .DO(ram16s_inst_781_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3127),
    .CLK(clk)
);

defparam ram16s_inst_781.INIT_0 = 16'h0000;
defparam ram16s_inst_781.INIT_1 = 16'h0000;
defparam ram16s_inst_781.INIT_2 = 16'h0000;
defparam ram16s_inst_781.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_782 (
    .DO(ram16s_inst_782_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3131),
    .CLK(clk)
);

defparam ram16s_inst_782.INIT_0 = 16'h0000;
defparam ram16s_inst_782.INIT_1 = 16'h0000;
defparam ram16s_inst_782.INIT_2 = 16'h0000;
defparam ram16s_inst_782.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_783 (
    .DO(ram16s_inst_783_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3135),
    .CLK(clk)
);

defparam ram16s_inst_783.INIT_0 = 16'h0000;
defparam ram16s_inst_783.INIT_1 = 16'h0000;
defparam ram16s_inst_783.INIT_2 = 16'h0000;
defparam ram16s_inst_783.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_784 (
    .DO(ram16s_inst_784_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3139),
    .CLK(clk)
);

defparam ram16s_inst_784.INIT_0 = 16'h0000;
defparam ram16s_inst_784.INIT_1 = 16'h0000;
defparam ram16s_inst_784.INIT_2 = 16'h0000;
defparam ram16s_inst_784.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_785 (
    .DO(ram16s_inst_785_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3143),
    .CLK(clk)
);

defparam ram16s_inst_785.INIT_0 = 16'h0000;
defparam ram16s_inst_785.INIT_1 = 16'h0000;
defparam ram16s_inst_785.INIT_2 = 16'h0000;
defparam ram16s_inst_785.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_786 (
    .DO(ram16s_inst_786_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3147),
    .CLK(clk)
);

defparam ram16s_inst_786.INIT_0 = 16'h0000;
defparam ram16s_inst_786.INIT_1 = 16'h0000;
defparam ram16s_inst_786.INIT_2 = 16'h0000;
defparam ram16s_inst_786.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_787 (
    .DO(ram16s_inst_787_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3151),
    .CLK(clk)
);

defparam ram16s_inst_787.INIT_0 = 16'h0000;
defparam ram16s_inst_787.INIT_1 = 16'h0000;
defparam ram16s_inst_787.INIT_2 = 16'h0000;
defparam ram16s_inst_787.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_788 (
    .DO(ram16s_inst_788_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3155),
    .CLK(clk)
);

defparam ram16s_inst_788.INIT_0 = 16'h0000;
defparam ram16s_inst_788.INIT_1 = 16'h0000;
defparam ram16s_inst_788.INIT_2 = 16'h0000;
defparam ram16s_inst_788.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_789 (
    .DO(ram16s_inst_789_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3159),
    .CLK(clk)
);

defparam ram16s_inst_789.INIT_0 = 16'h0000;
defparam ram16s_inst_789.INIT_1 = 16'h0000;
defparam ram16s_inst_789.INIT_2 = 16'h0000;
defparam ram16s_inst_789.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_790 (
    .DO(ram16s_inst_790_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3163),
    .CLK(clk)
);

defparam ram16s_inst_790.INIT_0 = 16'h0000;
defparam ram16s_inst_790.INIT_1 = 16'h0000;
defparam ram16s_inst_790.INIT_2 = 16'h0000;
defparam ram16s_inst_790.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_791 (
    .DO(ram16s_inst_791_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3167),
    .CLK(clk)
);

defparam ram16s_inst_791.INIT_0 = 16'h0000;
defparam ram16s_inst_791.INIT_1 = 16'h0000;
defparam ram16s_inst_791.INIT_2 = 16'h0000;
defparam ram16s_inst_791.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_792 (
    .DO(ram16s_inst_792_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3171),
    .CLK(clk)
);

defparam ram16s_inst_792.INIT_0 = 16'h0000;
defparam ram16s_inst_792.INIT_1 = 16'h0000;
defparam ram16s_inst_792.INIT_2 = 16'h0000;
defparam ram16s_inst_792.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_793 (
    .DO(ram16s_inst_793_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3175),
    .CLK(clk)
);

defparam ram16s_inst_793.INIT_0 = 16'h0000;
defparam ram16s_inst_793.INIT_1 = 16'h0000;
defparam ram16s_inst_793.INIT_2 = 16'h0000;
defparam ram16s_inst_793.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_794 (
    .DO(ram16s_inst_794_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3179),
    .CLK(clk)
);

defparam ram16s_inst_794.INIT_0 = 16'h0000;
defparam ram16s_inst_794.INIT_1 = 16'h0000;
defparam ram16s_inst_794.INIT_2 = 16'h0000;
defparam ram16s_inst_794.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_795 (
    .DO(ram16s_inst_795_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3183),
    .CLK(clk)
);

defparam ram16s_inst_795.INIT_0 = 16'h0000;
defparam ram16s_inst_795.INIT_1 = 16'h0000;
defparam ram16s_inst_795.INIT_2 = 16'h0000;
defparam ram16s_inst_795.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_796 (
    .DO(ram16s_inst_796_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3187),
    .CLK(clk)
);

defparam ram16s_inst_796.INIT_0 = 16'h0000;
defparam ram16s_inst_796.INIT_1 = 16'h0000;
defparam ram16s_inst_796.INIT_2 = 16'h0000;
defparam ram16s_inst_796.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_797 (
    .DO(ram16s_inst_797_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3191),
    .CLK(clk)
);

defparam ram16s_inst_797.INIT_0 = 16'h0000;
defparam ram16s_inst_797.INIT_1 = 16'h0000;
defparam ram16s_inst_797.INIT_2 = 16'h0000;
defparam ram16s_inst_797.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_798 (
    .DO(ram16s_inst_798_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3195),
    .CLK(clk)
);

defparam ram16s_inst_798.INIT_0 = 16'h0000;
defparam ram16s_inst_798.INIT_1 = 16'h0000;
defparam ram16s_inst_798.INIT_2 = 16'h0000;
defparam ram16s_inst_798.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_799 (
    .DO(ram16s_inst_799_dout[2:0]),
    .DI(di[2:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_3199),
    .CLK(clk)
);

defparam ram16s_inst_799.INIT_0 = 16'h0000;
defparam ram16s_inst_799.INIT_1 = 16'h0000;
defparam ram16s_inst_799.INIT_2 = 16'h0000;
defparam ram16s_inst_799.INIT_3 = 16'h0000;

MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(ram16s_inst_0_dout[0]),
  .I1(ram16s_inst_1_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(ram16s_inst_2_dout[0]),
  .I1(ram16s_inst_3_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(ram16s_inst_4_dout[0]),
  .I1(ram16s_inst_5_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(ram16s_inst_6_dout[0]),
  .I1(ram16s_inst_7_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(ram16s_inst_8_dout[0]),
  .I1(ram16s_inst_9_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(ram16s_inst_10_dout[0]),
  .I1(ram16s_inst_11_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(ram16s_inst_12_dout[0]),
  .I1(ram16s_inst_13_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(ram16s_inst_14_dout[0]),
  .I1(ram16s_inst_15_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(ram16s_inst_16_dout[0]),
  .I1(ram16s_inst_17_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(ram16s_inst_18_dout[0]),
  .I1(ram16s_inst_19_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(ram16s_inst_20_dout[0]),
  .I1(ram16s_inst_21_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(ram16s_inst_22_dout[0]),
  .I1(ram16s_inst_23_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(ram16s_inst_24_dout[0]),
  .I1(ram16s_inst_25_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(ram16s_inst_26_dout[0]),
  .I1(ram16s_inst_27_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(ram16s_inst_28_dout[0]),
  .I1(ram16s_inst_29_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(ram16s_inst_30_dout[0]),
  .I1(ram16s_inst_31_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(ram16s_inst_32_dout[0]),
  .I1(ram16s_inst_33_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(ram16s_inst_34_dout[0]),
  .I1(ram16s_inst_35_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(ram16s_inst_36_dout[0]),
  .I1(ram16s_inst_37_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(ram16s_inst_38_dout[0]),
  .I1(ram16s_inst_39_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(ram16s_inst_40_dout[0]),
  .I1(ram16s_inst_41_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(ram16s_inst_42_dout[0]),
  .I1(ram16s_inst_43_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(ram16s_inst_44_dout[0]),
  .I1(ram16s_inst_45_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(ram16s_inst_46_dout[0]),
  .I1(ram16s_inst_47_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(ram16s_inst_48_dout[0]),
  .I1(ram16s_inst_49_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(ram16s_inst_50_dout[0]),
  .I1(ram16s_inst_51_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(ram16s_inst_52_dout[0]),
  .I1(ram16s_inst_53_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(ram16s_inst_54_dout[0]),
  .I1(ram16s_inst_55_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(ram16s_inst_56_dout[0]),
  .I1(ram16s_inst_57_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(ram16s_inst_58_dout[0]),
  .I1(ram16s_inst_59_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(ram16s_inst_60_dout[0]),
  .I1(ram16s_inst_61_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(ram16s_inst_62_dout[0]),
  .I1(ram16s_inst_63_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(ram16s_inst_64_dout[0]),
  .I1(ram16s_inst_65_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(ram16s_inst_66_dout[0]),
  .I1(ram16s_inst_67_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(ram16s_inst_68_dout[0]),
  .I1(ram16s_inst_69_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(ram16s_inst_70_dout[0]),
  .I1(ram16s_inst_71_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(ram16s_inst_72_dout[0]),
  .I1(ram16s_inst_73_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(ram16s_inst_74_dout[0]),
  .I1(ram16s_inst_75_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(ram16s_inst_76_dout[0]),
  .I1(ram16s_inst_77_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(ram16s_inst_78_dout[0]),
  .I1(ram16s_inst_79_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(ram16s_inst_80_dout[0]),
  .I1(ram16s_inst_81_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(ram16s_inst_82_dout[0]),
  .I1(ram16s_inst_83_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(ram16s_inst_84_dout[0]),
  .I1(ram16s_inst_85_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(ram16s_inst_86_dout[0]),
  .I1(ram16s_inst_87_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(ram16s_inst_88_dout[0]),
  .I1(ram16s_inst_89_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(ram16s_inst_90_dout[0]),
  .I1(ram16s_inst_91_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(ram16s_inst_92_dout[0]),
  .I1(ram16s_inst_93_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(ram16s_inst_94_dout[0]),
  .I1(ram16s_inst_95_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(ram16s_inst_96_dout[0]),
  .I1(ram16s_inst_97_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(ram16s_inst_98_dout[0]),
  .I1(ram16s_inst_99_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(ram16s_inst_100_dout[0]),
  .I1(ram16s_inst_101_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(ram16s_inst_102_dout[0]),
  .I1(ram16s_inst_103_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(ram16s_inst_104_dout[0]),
  .I1(ram16s_inst_105_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(ram16s_inst_106_dout[0]),
  .I1(ram16s_inst_107_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(ram16s_inst_108_dout[0]),
  .I1(ram16s_inst_109_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(ram16s_inst_110_dout[0]),
  .I1(ram16s_inst_111_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(ram16s_inst_112_dout[0]),
  .I1(ram16s_inst_113_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(ram16s_inst_114_dout[0]),
  .I1(ram16s_inst_115_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(ram16s_inst_116_dout[0]),
  .I1(ram16s_inst_117_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(ram16s_inst_118_dout[0]),
  .I1(ram16s_inst_119_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(ram16s_inst_120_dout[0]),
  .I1(ram16s_inst_121_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(ram16s_inst_122_dout[0]),
  .I1(ram16s_inst_123_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(ram16s_inst_124_dout[0]),
  .I1(ram16s_inst_125_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(ram16s_inst_126_dout[0]),
  .I1(ram16s_inst_127_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(ram16s_inst_128_dout[0]),
  .I1(ram16s_inst_129_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(ram16s_inst_130_dout[0]),
  .I1(ram16s_inst_131_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(ram16s_inst_132_dout[0]),
  .I1(ram16s_inst_133_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(ram16s_inst_134_dout[0]),
  .I1(ram16s_inst_135_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(ram16s_inst_136_dout[0]),
  .I1(ram16s_inst_137_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(ram16s_inst_138_dout[0]),
  .I1(ram16s_inst_139_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(ram16s_inst_140_dout[0]),
  .I1(ram16s_inst_141_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(ram16s_inst_142_dout[0]),
  .I1(ram16s_inst_143_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(ram16s_inst_144_dout[0]),
  .I1(ram16s_inst_145_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(ram16s_inst_146_dout[0]),
  .I1(ram16s_inst_147_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(ram16s_inst_148_dout[0]),
  .I1(ram16s_inst_149_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(ram16s_inst_150_dout[0]),
  .I1(ram16s_inst_151_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(ram16s_inst_152_dout[0]),
  .I1(ram16s_inst_153_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(ram16s_inst_154_dout[0]),
  .I1(ram16s_inst_155_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(ram16s_inst_156_dout[0]),
  .I1(ram16s_inst_157_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(ram16s_inst_158_dout[0]),
  .I1(ram16s_inst_159_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(ram16s_inst_160_dout[0]),
  .I1(ram16s_inst_161_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(ram16s_inst_162_dout[0]),
  .I1(ram16s_inst_163_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(ram16s_inst_164_dout[0]),
  .I1(ram16s_inst_165_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(ram16s_inst_166_dout[0]),
  .I1(ram16s_inst_167_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(ram16s_inst_168_dout[0]),
  .I1(ram16s_inst_169_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(ram16s_inst_170_dout[0]),
  .I1(ram16s_inst_171_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(ram16s_inst_172_dout[0]),
  .I1(ram16s_inst_173_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(ram16s_inst_174_dout[0]),
  .I1(ram16s_inst_175_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(ram16s_inst_176_dout[0]),
  .I1(ram16s_inst_177_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(ram16s_inst_178_dout[0]),
  .I1(ram16s_inst_179_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(ram16s_inst_180_dout[0]),
  .I1(ram16s_inst_181_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(ram16s_inst_182_dout[0]),
  .I1(ram16s_inst_183_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(ram16s_inst_184_dout[0]),
  .I1(ram16s_inst_185_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(ram16s_inst_186_dout[0]),
  .I1(ram16s_inst_187_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(ram16s_inst_188_dout[0]),
  .I1(ram16s_inst_189_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(ram16s_inst_190_dout[0]),
  .I1(ram16s_inst_191_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(ram16s_inst_192_dout[0]),
  .I1(ram16s_inst_193_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(ram16s_inst_194_dout[0]),
  .I1(ram16s_inst_195_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(ram16s_inst_196_dout[0]),
  .I1(ram16s_inst_197_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(ram16s_inst_198_dout[0]),
  .I1(ram16s_inst_199_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(ram16s_inst_200_dout[0]),
  .I1(ram16s_inst_201_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(ram16s_inst_202_dout[0]),
  .I1(ram16s_inst_203_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(ram16s_inst_204_dout[0]),
  .I1(ram16s_inst_205_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(ram16s_inst_206_dout[0]),
  .I1(ram16s_inst_207_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_104 (
  .O(mux_o_104),
  .I0(ram16s_inst_208_dout[0]),
  .I1(ram16s_inst_209_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(ram16s_inst_210_dout[0]),
  .I1(ram16s_inst_211_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(ram16s_inst_212_dout[0]),
  .I1(ram16s_inst_213_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(ram16s_inst_214_dout[0]),
  .I1(ram16s_inst_215_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(ram16s_inst_216_dout[0]),
  .I1(ram16s_inst_217_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(ram16s_inst_218_dout[0]),
  .I1(ram16s_inst_219_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(ram16s_inst_220_dout[0]),
  .I1(ram16s_inst_221_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(ram16s_inst_222_dout[0]),
  .I1(ram16s_inst_223_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(ram16s_inst_224_dout[0]),
  .I1(ram16s_inst_225_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(ram16s_inst_226_dout[0]),
  .I1(ram16s_inst_227_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(ram16s_inst_228_dout[0]),
  .I1(ram16s_inst_229_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(ram16s_inst_230_dout[0]),
  .I1(ram16s_inst_231_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(ram16s_inst_232_dout[0]),
  .I1(ram16s_inst_233_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(ram16s_inst_234_dout[0]),
  .I1(ram16s_inst_235_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(ram16s_inst_236_dout[0]),
  .I1(ram16s_inst_237_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(ram16s_inst_238_dout[0]),
  .I1(ram16s_inst_239_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(ram16s_inst_240_dout[0]),
  .I1(ram16s_inst_241_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(ram16s_inst_242_dout[0]),
  .I1(ram16s_inst_243_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(ram16s_inst_244_dout[0]),
  .I1(ram16s_inst_245_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_123 (
  .O(mux_o_123),
  .I0(ram16s_inst_246_dout[0]),
  .I1(ram16s_inst_247_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(ram16s_inst_248_dout[0]),
  .I1(ram16s_inst_249_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_125 (
  .O(mux_o_125),
  .I0(ram16s_inst_250_dout[0]),
  .I1(ram16s_inst_251_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(ram16s_inst_252_dout[0]),
  .I1(ram16s_inst_253_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(ram16s_inst_254_dout[0]),
  .I1(ram16s_inst_255_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(ram16s_inst_256_dout[0]),
  .I1(ram16s_inst_257_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(ram16s_inst_258_dout[0]),
  .I1(ram16s_inst_259_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(ram16s_inst_260_dout[0]),
  .I1(ram16s_inst_261_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(ram16s_inst_262_dout[0]),
  .I1(ram16s_inst_263_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(ram16s_inst_264_dout[0]),
  .I1(ram16s_inst_265_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(ram16s_inst_266_dout[0]),
  .I1(ram16s_inst_267_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(ram16s_inst_268_dout[0]),
  .I1(ram16s_inst_269_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(ram16s_inst_270_dout[0]),
  .I1(ram16s_inst_271_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(ram16s_inst_272_dout[0]),
  .I1(ram16s_inst_273_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(ram16s_inst_274_dout[0]),
  .I1(ram16s_inst_275_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(ram16s_inst_276_dout[0]),
  .I1(ram16s_inst_277_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(ram16s_inst_278_dout[0]),
  .I1(ram16s_inst_279_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(ram16s_inst_280_dout[0]),
  .I1(ram16s_inst_281_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(ram16s_inst_282_dout[0]),
  .I1(ram16s_inst_283_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(ram16s_inst_284_dout[0]),
  .I1(ram16s_inst_285_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(ram16s_inst_286_dout[0]),
  .I1(ram16s_inst_287_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(ram16s_inst_288_dout[0]),
  .I1(ram16s_inst_289_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(ram16s_inst_290_dout[0]),
  .I1(ram16s_inst_291_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(ram16s_inst_292_dout[0]),
  .I1(ram16s_inst_293_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(ram16s_inst_294_dout[0]),
  .I1(ram16s_inst_295_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(ram16s_inst_296_dout[0]),
  .I1(ram16s_inst_297_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(ram16s_inst_298_dout[0]),
  .I1(ram16s_inst_299_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(ram16s_inst_300_dout[0]),
  .I1(ram16s_inst_301_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(ram16s_inst_302_dout[0]),
  .I1(ram16s_inst_303_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(ram16s_inst_304_dout[0]),
  .I1(ram16s_inst_305_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(ram16s_inst_306_dout[0]),
  .I1(ram16s_inst_307_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(ram16s_inst_308_dout[0]),
  .I1(ram16s_inst_309_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(ram16s_inst_310_dout[0]),
  .I1(ram16s_inst_311_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(ram16s_inst_312_dout[0]),
  .I1(ram16s_inst_313_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(ram16s_inst_314_dout[0]),
  .I1(ram16s_inst_315_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(ram16s_inst_316_dout[0]),
  .I1(ram16s_inst_317_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(ram16s_inst_318_dout[0]),
  .I1(ram16s_inst_319_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(ram16s_inst_320_dout[0]),
  .I1(ram16s_inst_321_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(ram16s_inst_322_dout[0]),
  .I1(ram16s_inst_323_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(ram16s_inst_324_dout[0]),
  .I1(ram16s_inst_325_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(ram16s_inst_326_dout[0]),
  .I1(ram16s_inst_327_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_164 (
  .O(mux_o_164),
  .I0(ram16s_inst_328_dout[0]),
  .I1(ram16s_inst_329_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(ram16s_inst_330_dout[0]),
  .I1(ram16s_inst_331_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(ram16s_inst_332_dout[0]),
  .I1(ram16s_inst_333_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(ram16s_inst_334_dout[0]),
  .I1(ram16s_inst_335_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(ram16s_inst_336_dout[0]),
  .I1(ram16s_inst_337_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(ram16s_inst_338_dout[0]),
  .I1(ram16s_inst_339_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(ram16s_inst_340_dout[0]),
  .I1(ram16s_inst_341_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(ram16s_inst_342_dout[0]),
  .I1(ram16s_inst_343_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(ram16s_inst_344_dout[0]),
  .I1(ram16s_inst_345_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(ram16s_inst_346_dout[0]),
  .I1(ram16s_inst_347_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(ram16s_inst_348_dout[0]),
  .I1(ram16s_inst_349_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(ram16s_inst_350_dout[0]),
  .I1(ram16s_inst_351_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(ram16s_inst_352_dout[0]),
  .I1(ram16s_inst_353_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(ram16s_inst_354_dout[0]),
  .I1(ram16s_inst_355_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(ram16s_inst_356_dout[0]),
  .I1(ram16s_inst_357_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(ram16s_inst_358_dout[0]),
  .I1(ram16s_inst_359_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(ram16s_inst_360_dout[0]),
  .I1(ram16s_inst_361_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(ram16s_inst_362_dout[0]),
  .I1(ram16s_inst_363_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(ram16s_inst_364_dout[0]),
  .I1(ram16s_inst_365_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(ram16s_inst_366_dout[0]),
  .I1(ram16s_inst_367_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(ram16s_inst_368_dout[0]),
  .I1(ram16s_inst_369_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(ram16s_inst_370_dout[0]),
  .I1(ram16s_inst_371_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(ram16s_inst_372_dout[0]),
  .I1(ram16s_inst_373_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(ram16s_inst_374_dout[0]),
  .I1(ram16s_inst_375_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(ram16s_inst_376_dout[0]),
  .I1(ram16s_inst_377_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(ram16s_inst_378_dout[0]),
  .I1(ram16s_inst_379_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(ram16s_inst_380_dout[0]),
  .I1(ram16s_inst_381_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(ram16s_inst_382_dout[0]),
  .I1(ram16s_inst_383_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(ram16s_inst_384_dout[0]),
  .I1(ram16s_inst_385_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(ram16s_inst_386_dout[0]),
  .I1(ram16s_inst_387_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(ram16s_inst_388_dout[0]),
  .I1(ram16s_inst_389_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(ram16s_inst_390_dout[0]),
  .I1(ram16s_inst_391_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(ram16s_inst_392_dout[0]),
  .I1(ram16s_inst_393_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(ram16s_inst_394_dout[0]),
  .I1(ram16s_inst_395_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(ram16s_inst_396_dout[0]),
  .I1(ram16s_inst_397_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(ram16s_inst_398_dout[0]),
  .I1(ram16s_inst_399_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(ram16s_inst_400_dout[0]),
  .I1(ram16s_inst_401_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(ram16s_inst_402_dout[0]),
  .I1(ram16s_inst_403_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(ram16s_inst_404_dout[0]),
  .I1(ram16s_inst_405_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(ram16s_inst_406_dout[0]),
  .I1(ram16s_inst_407_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(ram16s_inst_408_dout[0]),
  .I1(ram16s_inst_409_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(ram16s_inst_410_dout[0]),
  .I1(ram16s_inst_411_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(ram16s_inst_412_dout[0]),
  .I1(ram16s_inst_413_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(ram16s_inst_414_dout[0]),
  .I1(ram16s_inst_415_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(ram16s_inst_416_dout[0]),
  .I1(ram16s_inst_417_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_209 (
  .O(mux_o_209),
  .I0(ram16s_inst_418_dout[0]),
  .I1(ram16s_inst_419_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(ram16s_inst_420_dout[0]),
  .I1(ram16s_inst_421_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(ram16s_inst_422_dout[0]),
  .I1(ram16s_inst_423_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(ram16s_inst_424_dout[0]),
  .I1(ram16s_inst_425_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(ram16s_inst_426_dout[0]),
  .I1(ram16s_inst_427_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(ram16s_inst_428_dout[0]),
  .I1(ram16s_inst_429_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(ram16s_inst_430_dout[0]),
  .I1(ram16s_inst_431_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_216 (
  .O(mux_o_216),
  .I0(ram16s_inst_432_dout[0]),
  .I1(ram16s_inst_433_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(ram16s_inst_434_dout[0]),
  .I1(ram16s_inst_435_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(ram16s_inst_436_dout[0]),
  .I1(ram16s_inst_437_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(ram16s_inst_438_dout[0]),
  .I1(ram16s_inst_439_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(ram16s_inst_440_dout[0]),
  .I1(ram16s_inst_441_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(ram16s_inst_442_dout[0]),
  .I1(ram16s_inst_443_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(ram16s_inst_444_dout[0]),
  .I1(ram16s_inst_445_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(ram16s_inst_446_dout[0]),
  .I1(ram16s_inst_447_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_224 (
  .O(mux_o_224),
  .I0(ram16s_inst_448_dout[0]),
  .I1(ram16s_inst_449_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(ram16s_inst_450_dout[0]),
  .I1(ram16s_inst_451_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(ram16s_inst_452_dout[0]),
  .I1(ram16s_inst_453_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(ram16s_inst_454_dout[0]),
  .I1(ram16s_inst_455_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(ram16s_inst_456_dout[0]),
  .I1(ram16s_inst_457_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(ram16s_inst_458_dout[0]),
  .I1(ram16s_inst_459_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(ram16s_inst_460_dout[0]),
  .I1(ram16s_inst_461_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(ram16s_inst_462_dout[0]),
  .I1(ram16s_inst_463_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(ram16s_inst_464_dout[0]),
  .I1(ram16s_inst_465_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(ram16s_inst_466_dout[0]),
  .I1(ram16s_inst_467_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(ram16s_inst_468_dout[0]),
  .I1(ram16s_inst_469_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(ram16s_inst_470_dout[0]),
  .I1(ram16s_inst_471_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(ram16s_inst_472_dout[0]),
  .I1(ram16s_inst_473_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(ram16s_inst_474_dout[0]),
  .I1(ram16s_inst_475_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(ram16s_inst_476_dout[0]),
  .I1(ram16s_inst_477_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(ram16s_inst_478_dout[0]),
  .I1(ram16s_inst_479_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(ram16s_inst_480_dout[0]),
  .I1(ram16s_inst_481_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(ram16s_inst_482_dout[0]),
  .I1(ram16s_inst_483_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(ram16s_inst_484_dout[0]),
  .I1(ram16s_inst_485_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(ram16s_inst_486_dout[0]),
  .I1(ram16s_inst_487_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(ram16s_inst_488_dout[0]),
  .I1(ram16s_inst_489_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(ram16s_inst_490_dout[0]),
  .I1(ram16s_inst_491_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(ram16s_inst_492_dout[0]),
  .I1(ram16s_inst_493_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(ram16s_inst_494_dout[0]),
  .I1(ram16s_inst_495_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(ram16s_inst_496_dout[0]),
  .I1(ram16s_inst_497_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(ram16s_inst_498_dout[0]),
  .I1(ram16s_inst_499_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(ram16s_inst_500_dout[0]),
  .I1(ram16s_inst_501_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_251 (
  .O(mux_o_251),
  .I0(ram16s_inst_502_dout[0]),
  .I1(ram16s_inst_503_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(ram16s_inst_504_dout[0]),
  .I1(ram16s_inst_505_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(ram16s_inst_506_dout[0]),
  .I1(ram16s_inst_507_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_254 (
  .O(mux_o_254),
  .I0(ram16s_inst_508_dout[0]),
  .I1(ram16s_inst_509_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(ram16s_inst_510_dout[0]),
  .I1(ram16s_inst_511_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_256 (
  .O(mux_o_256),
  .I0(ram16s_inst_512_dout[0]),
  .I1(ram16s_inst_513_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(ram16s_inst_514_dout[0]),
  .I1(ram16s_inst_515_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(ram16s_inst_516_dout[0]),
  .I1(ram16s_inst_517_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(ram16s_inst_518_dout[0]),
  .I1(ram16s_inst_519_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(ram16s_inst_520_dout[0]),
  .I1(ram16s_inst_521_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(ram16s_inst_522_dout[0]),
  .I1(ram16s_inst_523_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_262 (
  .O(mux_o_262),
  .I0(ram16s_inst_524_dout[0]),
  .I1(ram16s_inst_525_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(ram16s_inst_526_dout[0]),
  .I1(ram16s_inst_527_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(ram16s_inst_528_dout[0]),
  .I1(ram16s_inst_529_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_265 (
  .O(mux_o_265),
  .I0(ram16s_inst_530_dout[0]),
  .I1(ram16s_inst_531_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(ram16s_inst_532_dout[0]),
  .I1(ram16s_inst_533_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(ram16s_inst_534_dout[0]),
  .I1(ram16s_inst_535_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(ram16s_inst_536_dout[0]),
  .I1(ram16s_inst_537_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_269 (
  .O(mux_o_269),
  .I0(ram16s_inst_538_dout[0]),
  .I1(ram16s_inst_539_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(ram16s_inst_540_dout[0]),
  .I1(ram16s_inst_541_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(ram16s_inst_542_dout[0]),
  .I1(ram16s_inst_543_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_272 (
  .O(mux_o_272),
  .I0(ram16s_inst_544_dout[0]),
  .I1(ram16s_inst_545_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(ram16s_inst_546_dout[0]),
  .I1(ram16s_inst_547_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(ram16s_inst_548_dout[0]),
  .I1(ram16s_inst_549_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(ram16s_inst_550_dout[0]),
  .I1(ram16s_inst_551_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_276 (
  .O(mux_o_276),
  .I0(ram16s_inst_552_dout[0]),
  .I1(ram16s_inst_553_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(ram16s_inst_554_dout[0]),
  .I1(ram16s_inst_555_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_278 (
  .O(mux_o_278),
  .I0(ram16s_inst_556_dout[0]),
  .I1(ram16s_inst_557_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_279 (
  .O(mux_o_279),
  .I0(ram16s_inst_558_dout[0]),
  .I1(ram16s_inst_559_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(ram16s_inst_560_dout[0]),
  .I1(ram16s_inst_561_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(ram16s_inst_562_dout[0]),
  .I1(ram16s_inst_563_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(ram16s_inst_564_dout[0]),
  .I1(ram16s_inst_565_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(ram16s_inst_566_dout[0]),
  .I1(ram16s_inst_567_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_284 (
  .O(mux_o_284),
  .I0(ram16s_inst_568_dout[0]),
  .I1(ram16s_inst_569_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(ram16s_inst_570_dout[0]),
  .I1(ram16s_inst_571_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(ram16s_inst_572_dout[0]),
  .I1(ram16s_inst_573_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(ram16s_inst_574_dout[0]),
  .I1(ram16s_inst_575_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(ram16s_inst_576_dout[0]),
  .I1(ram16s_inst_577_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(ram16s_inst_578_dout[0]),
  .I1(ram16s_inst_579_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(ram16s_inst_580_dout[0]),
  .I1(ram16s_inst_581_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(ram16s_inst_582_dout[0]),
  .I1(ram16s_inst_583_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(ram16s_inst_584_dout[0]),
  .I1(ram16s_inst_585_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_293 (
  .O(mux_o_293),
  .I0(ram16s_inst_586_dout[0]),
  .I1(ram16s_inst_587_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(ram16s_inst_588_dout[0]),
  .I1(ram16s_inst_589_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(ram16s_inst_590_dout[0]),
  .I1(ram16s_inst_591_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(ram16s_inst_592_dout[0]),
  .I1(ram16s_inst_593_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(ram16s_inst_594_dout[0]),
  .I1(ram16s_inst_595_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(ram16s_inst_596_dout[0]),
  .I1(ram16s_inst_597_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(ram16s_inst_598_dout[0]),
  .I1(ram16s_inst_599_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(ram16s_inst_600_dout[0]),
  .I1(ram16s_inst_601_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(ram16s_inst_602_dout[0]),
  .I1(ram16s_inst_603_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(ram16s_inst_604_dout[0]),
  .I1(ram16s_inst_605_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(ram16s_inst_606_dout[0]),
  .I1(ram16s_inst_607_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_304 (
  .O(mux_o_304),
  .I0(ram16s_inst_608_dout[0]),
  .I1(ram16s_inst_609_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(ram16s_inst_610_dout[0]),
  .I1(ram16s_inst_611_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(ram16s_inst_612_dout[0]),
  .I1(ram16s_inst_613_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(ram16s_inst_614_dout[0]),
  .I1(ram16s_inst_615_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(ram16s_inst_616_dout[0]),
  .I1(ram16s_inst_617_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(ram16s_inst_618_dout[0]),
  .I1(ram16s_inst_619_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(ram16s_inst_620_dout[0]),
  .I1(ram16s_inst_621_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(ram16s_inst_622_dout[0]),
  .I1(ram16s_inst_623_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(ram16s_inst_624_dout[0]),
  .I1(ram16s_inst_625_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(ram16s_inst_626_dout[0]),
  .I1(ram16s_inst_627_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_314 (
  .O(mux_o_314),
  .I0(ram16s_inst_628_dout[0]),
  .I1(ram16s_inst_629_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(ram16s_inst_630_dout[0]),
  .I1(ram16s_inst_631_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(ram16s_inst_632_dout[0]),
  .I1(ram16s_inst_633_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(ram16s_inst_634_dout[0]),
  .I1(ram16s_inst_635_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(ram16s_inst_636_dout[0]),
  .I1(ram16s_inst_637_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(ram16s_inst_638_dout[0]),
  .I1(ram16s_inst_639_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(ram16s_inst_640_dout[0]),
  .I1(ram16s_inst_641_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_321 (
  .O(mux_o_321),
  .I0(ram16s_inst_642_dout[0]),
  .I1(ram16s_inst_643_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(ram16s_inst_644_dout[0]),
  .I1(ram16s_inst_645_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(ram16s_inst_646_dout[0]),
  .I1(ram16s_inst_647_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(ram16s_inst_648_dout[0]),
  .I1(ram16s_inst_649_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(ram16s_inst_650_dout[0]),
  .I1(ram16s_inst_651_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(ram16s_inst_652_dout[0]),
  .I1(ram16s_inst_653_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(ram16s_inst_654_dout[0]),
  .I1(ram16s_inst_655_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_328 (
  .O(mux_o_328),
  .I0(ram16s_inst_656_dout[0]),
  .I1(ram16s_inst_657_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_329 (
  .O(mux_o_329),
  .I0(ram16s_inst_658_dout[0]),
  .I1(ram16s_inst_659_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(ram16s_inst_660_dout[0]),
  .I1(ram16s_inst_661_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(ram16s_inst_662_dout[0]),
  .I1(ram16s_inst_663_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(ram16s_inst_664_dout[0]),
  .I1(ram16s_inst_665_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(ram16s_inst_666_dout[0]),
  .I1(ram16s_inst_667_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(ram16s_inst_668_dout[0]),
  .I1(ram16s_inst_669_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_335 (
  .O(mux_o_335),
  .I0(ram16s_inst_670_dout[0]),
  .I1(ram16s_inst_671_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(ram16s_inst_672_dout[0]),
  .I1(ram16s_inst_673_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(ram16s_inst_674_dout[0]),
  .I1(ram16s_inst_675_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(ram16s_inst_676_dout[0]),
  .I1(ram16s_inst_677_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(ram16s_inst_678_dout[0]),
  .I1(ram16s_inst_679_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(ram16s_inst_680_dout[0]),
  .I1(ram16s_inst_681_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(ram16s_inst_682_dout[0]),
  .I1(ram16s_inst_683_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(ram16s_inst_684_dout[0]),
  .I1(ram16s_inst_685_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(ram16s_inst_686_dout[0]),
  .I1(ram16s_inst_687_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(ram16s_inst_688_dout[0]),
  .I1(ram16s_inst_689_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(ram16s_inst_690_dout[0]),
  .I1(ram16s_inst_691_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(ram16s_inst_692_dout[0]),
  .I1(ram16s_inst_693_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(ram16s_inst_694_dout[0]),
  .I1(ram16s_inst_695_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(ram16s_inst_696_dout[0]),
  .I1(ram16s_inst_697_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_349 (
  .O(mux_o_349),
  .I0(ram16s_inst_698_dout[0]),
  .I1(ram16s_inst_699_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(ram16s_inst_700_dout[0]),
  .I1(ram16s_inst_701_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(ram16s_inst_702_dout[0]),
  .I1(ram16s_inst_703_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(ram16s_inst_704_dout[0]),
  .I1(ram16s_inst_705_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(ram16s_inst_706_dout[0]),
  .I1(ram16s_inst_707_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(ram16s_inst_708_dout[0]),
  .I1(ram16s_inst_709_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(ram16s_inst_710_dout[0]),
  .I1(ram16s_inst_711_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_356 (
  .O(mux_o_356),
  .I0(ram16s_inst_712_dout[0]),
  .I1(ram16s_inst_713_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(ram16s_inst_714_dout[0]),
  .I1(ram16s_inst_715_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(ram16s_inst_716_dout[0]),
  .I1(ram16s_inst_717_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(ram16s_inst_718_dout[0]),
  .I1(ram16s_inst_719_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(ram16s_inst_720_dout[0]),
  .I1(ram16s_inst_721_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(ram16s_inst_722_dout[0]),
  .I1(ram16s_inst_723_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(ram16s_inst_724_dout[0]),
  .I1(ram16s_inst_725_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_363 (
  .O(mux_o_363),
  .I0(ram16s_inst_726_dout[0]),
  .I1(ram16s_inst_727_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(ram16s_inst_728_dout[0]),
  .I1(ram16s_inst_729_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(ram16s_inst_730_dout[0]),
  .I1(ram16s_inst_731_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(ram16s_inst_732_dout[0]),
  .I1(ram16s_inst_733_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(ram16s_inst_734_dout[0]),
  .I1(ram16s_inst_735_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(ram16s_inst_736_dout[0]),
  .I1(ram16s_inst_737_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(ram16s_inst_738_dout[0]),
  .I1(ram16s_inst_739_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_370 (
  .O(mux_o_370),
  .I0(ram16s_inst_740_dout[0]),
  .I1(ram16s_inst_741_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_371 (
  .O(mux_o_371),
  .I0(ram16s_inst_742_dout[0]),
  .I1(ram16s_inst_743_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(ram16s_inst_744_dout[0]),
  .I1(ram16s_inst_745_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(ram16s_inst_746_dout[0]),
  .I1(ram16s_inst_747_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_374 (
  .O(mux_o_374),
  .I0(ram16s_inst_748_dout[0]),
  .I1(ram16s_inst_749_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(ram16s_inst_750_dout[0]),
  .I1(ram16s_inst_751_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(ram16s_inst_752_dout[0]),
  .I1(ram16s_inst_753_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_377 (
  .O(mux_o_377),
  .I0(ram16s_inst_754_dout[0]),
  .I1(ram16s_inst_755_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_378 (
  .O(mux_o_378),
  .I0(ram16s_inst_756_dout[0]),
  .I1(ram16s_inst_757_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_379 (
  .O(mux_o_379),
  .I0(ram16s_inst_758_dout[0]),
  .I1(ram16s_inst_759_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_380 (
  .O(mux_o_380),
  .I0(ram16s_inst_760_dout[0]),
  .I1(ram16s_inst_761_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_381 (
  .O(mux_o_381),
  .I0(ram16s_inst_762_dout[0]),
  .I1(ram16s_inst_763_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_382 (
  .O(mux_o_382),
  .I0(ram16s_inst_764_dout[0]),
  .I1(ram16s_inst_765_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_383 (
  .O(mux_o_383),
  .I0(ram16s_inst_766_dout[0]),
  .I1(ram16s_inst_767_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_384 (
  .O(mux_o_384),
  .I0(ram16s_inst_768_dout[0]),
  .I1(ram16s_inst_769_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_385 (
  .O(mux_o_385),
  .I0(ram16s_inst_770_dout[0]),
  .I1(ram16s_inst_771_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_386 (
  .O(mux_o_386),
  .I0(ram16s_inst_772_dout[0]),
  .I1(ram16s_inst_773_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_387 (
  .O(mux_o_387),
  .I0(ram16s_inst_774_dout[0]),
  .I1(ram16s_inst_775_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_388 (
  .O(mux_o_388),
  .I0(ram16s_inst_776_dout[0]),
  .I1(ram16s_inst_777_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_389 (
  .O(mux_o_389),
  .I0(ram16s_inst_778_dout[0]),
  .I1(ram16s_inst_779_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(ram16s_inst_780_dout[0]),
  .I1(ram16s_inst_781_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_391 (
  .O(mux_o_391),
  .I0(ram16s_inst_782_dout[0]),
  .I1(ram16s_inst_783_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(ram16s_inst_784_dout[0]),
  .I1(ram16s_inst_785_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(ram16s_inst_786_dout[0]),
  .I1(ram16s_inst_787_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(ram16s_inst_788_dout[0]),
  .I1(ram16s_inst_789_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(ram16s_inst_790_dout[0]),
  .I1(ram16s_inst_791_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(ram16s_inst_792_dout[0]),
  .I1(ram16s_inst_793_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(ram16s_inst_794_dout[0]),
  .I1(ram16s_inst_795_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_398 (
  .O(mux_o_398),
  .I0(ram16s_inst_796_dout[0]),
  .I1(ram16s_inst_797_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(ram16s_inst_798_dout[0]),
  .I1(ram16s_inst_799_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(ad[5])
);
MUX2 mux_inst_401 (
  .O(mux_o_401),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(ad[5])
);
MUX2 mux_inst_402 (
  .O(mux_o_402),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(ad[5])
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(ad[5])
);
MUX2 mux_inst_404 (
  .O(mux_o_404),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(ad[5])
);
MUX2 mux_inst_405 (
  .O(mux_o_405),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(ad[5])
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(ad[5])
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(ad[5])
);
MUX2 mux_inst_408 (
  .O(mux_o_408),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(ad[5])
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(ad[5])
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(mux_o_20),
  .I1(mux_o_21),
  .S0(ad[5])
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(mux_o_22),
  .I1(mux_o_23),
  .S0(ad[5])
);
MUX2 mux_inst_412 (
  .O(mux_o_412),
  .I0(mux_o_24),
  .I1(mux_o_25),
  .S0(ad[5])
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(mux_o_26),
  .I1(mux_o_27),
  .S0(ad[5])
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(mux_o_28),
  .I1(mux_o_29),
  .S0(ad[5])
);
MUX2 mux_inst_415 (
  .O(mux_o_415),
  .I0(mux_o_30),
  .I1(mux_o_31),
  .S0(ad[5])
);
MUX2 mux_inst_416 (
  .O(mux_o_416),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(ad[5])
);
MUX2 mux_inst_417 (
  .O(mux_o_417),
  .I0(mux_o_34),
  .I1(mux_o_35),
  .S0(ad[5])
);
MUX2 mux_inst_418 (
  .O(mux_o_418),
  .I0(mux_o_36),
  .I1(mux_o_37),
  .S0(ad[5])
);
MUX2 mux_inst_419 (
  .O(mux_o_419),
  .I0(mux_o_38),
  .I1(mux_o_39),
  .S0(ad[5])
);
MUX2 mux_inst_420 (
  .O(mux_o_420),
  .I0(mux_o_40),
  .I1(mux_o_41),
  .S0(ad[5])
);
MUX2 mux_inst_421 (
  .O(mux_o_421),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(ad[5])
);
MUX2 mux_inst_422 (
  .O(mux_o_422),
  .I0(mux_o_44),
  .I1(mux_o_45),
  .S0(ad[5])
);
MUX2 mux_inst_423 (
  .O(mux_o_423),
  .I0(mux_o_46),
  .I1(mux_o_47),
  .S0(ad[5])
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(mux_o_48),
  .I1(mux_o_49),
  .S0(ad[5])
);
MUX2 mux_inst_425 (
  .O(mux_o_425),
  .I0(mux_o_50),
  .I1(mux_o_51),
  .S0(ad[5])
);
MUX2 mux_inst_426 (
  .O(mux_o_426),
  .I0(mux_o_52),
  .I1(mux_o_53),
  .S0(ad[5])
);
MUX2 mux_inst_427 (
  .O(mux_o_427),
  .I0(mux_o_54),
  .I1(mux_o_55),
  .S0(ad[5])
);
MUX2 mux_inst_428 (
  .O(mux_o_428),
  .I0(mux_o_56),
  .I1(mux_o_57),
  .S0(ad[5])
);
MUX2 mux_inst_429 (
  .O(mux_o_429),
  .I0(mux_o_58),
  .I1(mux_o_59),
  .S0(ad[5])
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(ad[5])
);
MUX2 mux_inst_431 (
  .O(mux_o_431),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(ad[5])
);
MUX2 mux_inst_432 (
  .O(mux_o_432),
  .I0(mux_o_64),
  .I1(mux_o_65),
  .S0(ad[5])
);
MUX2 mux_inst_433 (
  .O(mux_o_433),
  .I0(mux_o_66),
  .I1(mux_o_67),
  .S0(ad[5])
);
MUX2 mux_inst_434 (
  .O(mux_o_434),
  .I0(mux_o_68),
  .I1(mux_o_69),
  .S0(ad[5])
);
MUX2 mux_inst_435 (
  .O(mux_o_435),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(ad[5])
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(ad[5])
);
MUX2 mux_inst_437 (
  .O(mux_o_437),
  .I0(mux_o_74),
  .I1(mux_o_75),
  .S0(ad[5])
);
MUX2 mux_inst_438 (
  .O(mux_o_438),
  .I0(mux_o_76),
  .I1(mux_o_77),
  .S0(ad[5])
);
MUX2 mux_inst_439 (
  .O(mux_o_439),
  .I0(mux_o_78),
  .I1(mux_o_79),
  .S0(ad[5])
);
MUX2 mux_inst_440 (
  .O(mux_o_440),
  .I0(mux_o_80),
  .I1(mux_o_81),
  .S0(ad[5])
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(mux_o_82),
  .I1(mux_o_83),
  .S0(ad[5])
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(mux_o_84),
  .I1(mux_o_85),
  .S0(ad[5])
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(mux_o_86),
  .I1(mux_o_87),
  .S0(ad[5])
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(mux_o_88),
  .I1(mux_o_89),
  .S0(ad[5])
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(ad[5])
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(mux_o_92),
  .I1(mux_o_93),
  .S0(ad[5])
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(mux_o_94),
  .I1(mux_o_95),
  .S0(ad[5])
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(mux_o_96),
  .I1(mux_o_97),
  .S0(ad[5])
);
MUX2 mux_inst_449 (
  .O(mux_o_449),
  .I0(mux_o_98),
  .I1(mux_o_99),
  .S0(ad[5])
);
MUX2 mux_inst_450 (
  .O(mux_o_450),
  .I0(mux_o_100),
  .I1(mux_o_101),
  .S0(ad[5])
);
MUX2 mux_inst_451 (
  .O(mux_o_451),
  .I0(mux_o_102),
  .I1(mux_o_103),
  .S0(ad[5])
);
MUX2 mux_inst_452 (
  .O(mux_o_452),
  .I0(mux_o_104),
  .I1(mux_o_105),
  .S0(ad[5])
);
MUX2 mux_inst_453 (
  .O(mux_o_453),
  .I0(mux_o_106),
  .I1(mux_o_107),
  .S0(ad[5])
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(mux_o_108),
  .I1(mux_o_109),
  .S0(ad[5])
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(mux_o_110),
  .I1(mux_o_111),
  .S0(ad[5])
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(mux_o_112),
  .I1(mux_o_113),
  .S0(ad[5])
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(mux_o_114),
  .I1(mux_o_115),
  .S0(ad[5])
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(mux_o_116),
  .I1(mux_o_117),
  .S0(ad[5])
);
MUX2 mux_inst_459 (
  .O(mux_o_459),
  .I0(mux_o_118),
  .I1(mux_o_119),
  .S0(ad[5])
);
MUX2 mux_inst_460 (
  .O(mux_o_460),
  .I0(mux_o_120),
  .I1(mux_o_121),
  .S0(ad[5])
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(mux_o_122),
  .I1(mux_o_123),
  .S0(ad[5])
);
MUX2 mux_inst_462 (
  .O(mux_o_462),
  .I0(mux_o_124),
  .I1(mux_o_125),
  .S0(ad[5])
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(ad[5])
);
MUX2 mux_inst_464 (
  .O(mux_o_464),
  .I0(mux_o_128),
  .I1(mux_o_129),
  .S0(ad[5])
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(ad[5])
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(mux_o_132),
  .I1(mux_o_133),
  .S0(ad[5])
);
MUX2 mux_inst_467 (
  .O(mux_o_467),
  .I0(mux_o_134),
  .I1(mux_o_135),
  .S0(ad[5])
);
MUX2 mux_inst_468 (
  .O(mux_o_468),
  .I0(mux_o_136),
  .I1(mux_o_137),
  .S0(ad[5])
);
MUX2 mux_inst_469 (
  .O(mux_o_469),
  .I0(mux_o_138),
  .I1(mux_o_139),
  .S0(ad[5])
);
MUX2 mux_inst_470 (
  .O(mux_o_470),
  .I0(mux_o_140),
  .I1(mux_o_141),
  .S0(ad[5])
);
MUX2 mux_inst_471 (
  .O(mux_o_471),
  .I0(mux_o_142),
  .I1(mux_o_143),
  .S0(ad[5])
);
MUX2 mux_inst_472 (
  .O(mux_o_472),
  .I0(mux_o_144),
  .I1(mux_o_145),
  .S0(ad[5])
);
MUX2 mux_inst_473 (
  .O(mux_o_473),
  .I0(mux_o_146),
  .I1(mux_o_147),
  .S0(ad[5])
);
MUX2 mux_inst_474 (
  .O(mux_o_474),
  .I0(mux_o_148),
  .I1(mux_o_149),
  .S0(ad[5])
);
MUX2 mux_inst_475 (
  .O(mux_o_475),
  .I0(mux_o_150),
  .I1(mux_o_151),
  .S0(ad[5])
);
MUX2 mux_inst_476 (
  .O(mux_o_476),
  .I0(mux_o_152),
  .I1(mux_o_153),
  .S0(ad[5])
);
MUX2 mux_inst_477 (
  .O(mux_o_477),
  .I0(mux_o_154),
  .I1(mux_o_155),
  .S0(ad[5])
);
MUX2 mux_inst_478 (
  .O(mux_o_478),
  .I0(mux_o_156),
  .I1(mux_o_157),
  .S0(ad[5])
);
MUX2 mux_inst_479 (
  .O(mux_o_479),
  .I0(mux_o_158),
  .I1(mux_o_159),
  .S0(ad[5])
);
MUX2 mux_inst_480 (
  .O(mux_o_480),
  .I0(mux_o_160),
  .I1(mux_o_161),
  .S0(ad[5])
);
MUX2 mux_inst_481 (
  .O(mux_o_481),
  .I0(mux_o_162),
  .I1(mux_o_163),
  .S0(ad[5])
);
MUX2 mux_inst_482 (
  .O(mux_o_482),
  .I0(mux_o_164),
  .I1(mux_o_165),
  .S0(ad[5])
);
MUX2 mux_inst_483 (
  .O(mux_o_483),
  .I0(mux_o_166),
  .I1(mux_o_167),
  .S0(ad[5])
);
MUX2 mux_inst_484 (
  .O(mux_o_484),
  .I0(mux_o_168),
  .I1(mux_o_169),
  .S0(ad[5])
);
MUX2 mux_inst_485 (
  .O(mux_o_485),
  .I0(mux_o_170),
  .I1(mux_o_171),
  .S0(ad[5])
);
MUX2 mux_inst_486 (
  .O(mux_o_486),
  .I0(mux_o_172),
  .I1(mux_o_173),
  .S0(ad[5])
);
MUX2 mux_inst_487 (
  .O(mux_o_487),
  .I0(mux_o_174),
  .I1(mux_o_175),
  .S0(ad[5])
);
MUX2 mux_inst_488 (
  .O(mux_o_488),
  .I0(mux_o_176),
  .I1(mux_o_177),
  .S0(ad[5])
);
MUX2 mux_inst_489 (
  .O(mux_o_489),
  .I0(mux_o_178),
  .I1(mux_o_179),
  .S0(ad[5])
);
MUX2 mux_inst_490 (
  .O(mux_o_490),
  .I0(mux_o_180),
  .I1(mux_o_181),
  .S0(ad[5])
);
MUX2 mux_inst_491 (
  .O(mux_o_491),
  .I0(mux_o_182),
  .I1(mux_o_183),
  .S0(ad[5])
);
MUX2 mux_inst_492 (
  .O(mux_o_492),
  .I0(mux_o_184),
  .I1(mux_o_185),
  .S0(ad[5])
);
MUX2 mux_inst_493 (
  .O(mux_o_493),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(ad[5])
);
MUX2 mux_inst_494 (
  .O(mux_o_494),
  .I0(mux_o_188),
  .I1(mux_o_189),
  .S0(ad[5])
);
MUX2 mux_inst_495 (
  .O(mux_o_495),
  .I0(mux_o_190),
  .I1(mux_o_191),
  .S0(ad[5])
);
MUX2 mux_inst_496 (
  .O(mux_o_496),
  .I0(mux_o_192),
  .I1(mux_o_193),
  .S0(ad[5])
);
MUX2 mux_inst_497 (
  .O(mux_o_497),
  .I0(mux_o_194),
  .I1(mux_o_195),
  .S0(ad[5])
);
MUX2 mux_inst_498 (
  .O(mux_o_498),
  .I0(mux_o_196),
  .I1(mux_o_197),
  .S0(ad[5])
);
MUX2 mux_inst_499 (
  .O(mux_o_499),
  .I0(mux_o_198),
  .I1(mux_o_199),
  .S0(ad[5])
);
MUX2 mux_inst_500 (
  .O(mux_o_500),
  .I0(mux_o_200),
  .I1(mux_o_201),
  .S0(ad[5])
);
MUX2 mux_inst_501 (
  .O(mux_o_501),
  .I0(mux_o_202),
  .I1(mux_o_203),
  .S0(ad[5])
);
MUX2 mux_inst_502 (
  .O(mux_o_502),
  .I0(mux_o_204),
  .I1(mux_o_205),
  .S0(ad[5])
);
MUX2 mux_inst_503 (
  .O(mux_o_503),
  .I0(mux_o_206),
  .I1(mux_o_207),
  .S0(ad[5])
);
MUX2 mux_inst_504 (
  .O(mux_o_504),
  .I0(mux_o_208),
  .I1(mux_o_209),
  .S0(ad[5])
);
MUX2 mux_inst_505 (
  .O(mux_o_505),
  .I0(mux_o_210),
  .I1(mux_o_211),
  .S0(ad[5])
);
MUX2 mux_inst_506 (
  .O(mux_o_506),
  .I0(mux_o_212),
  .I1(mux_o_213),
  .S0(ad[5])
);
MUX2 mux_inst_507 (
  .O(mux_o_507),
  .I0(mux_o_214),
  .I1(mux_o_215),
  .S0(ad[5])
);
MUX2 mux_inst_508 (
  .O(mux_o_508),
  .I0(mux_o_216),
  .I1(mux_o_217),
  .S0(ad[5])
);
MUX2 mux_inst_509 (
  .O(mux_o_509),
  .I0(mux_o_218),
  .I1(mux_o_219),
  .S0(ad[5])
);
MUX2 mux_inst_510 (
  .O(mux_o_510),
  .I0(mux_o_220),
  .I1(mux_o_221),
  .S0(ad[5])
);
MUX2 mux_inst_511 (
  .O(mux_o_511),
  .I0(mux_o_222),
  .I1(mux_o_223),
  .S0(ad[5])
);
MUX2 mux_inst_512 (
  .O(mux_o_512),
  .I0(mux_o_224),
  .I1(mux_o_225),
  .S0(ad[5])
);
MUX2 mux_inst_513 (
  .O(mux_o_513),
  .I0(mux_o_226),
  .I1(mux_o_227),
  .S0(ad[5])
);
MUX2 mux_inst_514 (
  .O(mux_o_514),
  .I0(mux_o_228),
  .I1(mux_o_229),
  .S0(ad[5])
);
MUX2 mux_inst_515 (
  .O(mux_o_515),
  .I0(mux_o_230),
  .I1(mux_o_231),
  .S0(ad[5])
);
MUX2 mux_inst_516 (
  .O(mux_o_516),
  .I0(mux_o_232),
  .I1(mux_o_233),
  .S0(ad[5])
);
MUX2 mux_inst_517 (
  .O(mux_o_517),
  .I0(mux_o_234),
  .I1(mux_o_235),
  .S0(ad[5])
);
MUX2 mux_inst_518 (
  .O(mux_o_518),
  .I0(mux_o_236),
  .I1(mux_o_237),
  .S0(ad[5])
);
MUX2 mux_inst_519 (
  .O(mux_o_519),
  .I0(mux_o_238),
  .I1(mux_o_239),
  .S0(ad[5])
);
MUX2 mux_inst_520 (
  .O(mux_o_520),
  .I0(mux_o_240),
  .I1(mux_o_241),
  .S0(ad[5])
);
MUX2 mux_inst_521 (
  .O(mux_o_521),
  .I0(mux_o_242),
  .I1(mux_o_243),
  .S0(ad[5])
);
MUX2 mux_inst_522 (
  .O(mux_o_522),
  .I0(mux_o_244),
  .I1(mux_o_245),
  .S0(ad[5])
);
MUX2 mux_inst_523 (
  .O(mux_o_523),
  .I0(mux_o_246),
  .I1(mux_o_247),
  .S0(ad[5])
);
MUX2 mux_inst_524 (
  .O(mux_o_524),
  .I0(mux_o_248),
  .I1(mux_o_249),
  .S0(ad[5])
);
MUX2 mux_inst_525 (
  .O(mux_o_525),
  .I0(mux_o_250),
  .I1(mux_o_251),
  .S0(ad[5])
);
MUX2 mux_inst_526 (
  .O(mux_o_526),
  .I0(mux_o_252),
  .I1(mux_o_253),
  .S0(ad[5])
);
MUX2 mux_inst_527 (
  .O(mux_o_527),
  .I0(mux_o_254),
  .I1(mux_o_255),
  .S0(ad[5])
);
MUX2 mux_inst_528 (
  .O(mux_o_528),
  .I0(mux_o_256),
  .I1(mux_o_257),
  .S0(ad[5])
);
MUX2 mux_inst_529 (
  .O(mux_o_529),
  .I0(mux_o_258),
  .I1(mux_o_259),
  .S0(ad[5])
);
MUX2 mux_inst_530 (
  .O(mux_o_530),
  .I0(mux_o_260),
  .I1(mux_o_261),
  .S0(ad[5])
);
MUX2 mux_inst_531 (
  .O(mux_o_531),
  .I0(mux_o_262),
  .I1(mux_o_263),
  .S0(ad[5])
);
MUX2 mux_inst_532 (
  .O(mux_o_532),
  .I0(mux_o_264),
  .I1(mux_o_265),
  .S0(ad[5])
);
MUX2 mux_inst_533 (
  .O(mux_o_533),
  .I0(mux_o_266),
  .I1(mux_o_267),
  .S0(ad[5])
);
MUX2 mux_inst_534 (
  .O(mux_o_534),
  .I0(mux_o_268),
  .I1(mux_o_269),
  .S0(ad[5])
);
MUX2 mux_inst_535 (
  .O(mux_o_535),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(ad[5])
);
MUX2 mux_inst_536 (
  .O(mux_o_536),
  .I0(mux_o_272),
  .I1(mux_o_273),
  .S0(ad[5])
);
MUX2 mux_inst_537 (
  .O(mux_o_537),
  .I0(mux_o_274),
  .I1(mux_o_275),
  .S0(ad[5])
);
MUX2 mux_inst_538 (
  .O(mux_o_538),
  .I0(mux_o_276),
  .I1(mux_o_277),
  .S0(ad[5])
);
MUX2 mux_inst_539 (
  .O(mux_o_539),
  .I0(mux_o_278),
  .I1(mux_o_279),
  .S0(ad[5])
);
MUX2 mux_inst_540 (
  .O(mux_o_540),
  .I0(mux_o_280),
  .I1(mux_o_281),
  .S0(ad[5])
);
MUX2 mux_inst_541 (
  .O(mux_o_541),
  .I0(mux_o_282),
  .I1(mux_o_283),
  .S0(ad[5])
);
MUX2 mux_inst_542 (
  .O(mux_o_542),
  .I0(mux_o_284),
  .I1(mux_o_285),
  .S0(ad[5])
);
MUX2 mux_inst_543 (
  .O(mux_o_543),
  .I0(mux_o_286),
  .I1(mux_o_287),
  .S0(ad[5])
);
MUX2 mux_inst_544 (
  .O(mux_o_544),
  .I0(mux_o_288),
  .I1(mux_o_289),
  .S0(ad[5])
);
MUX2 mux_inst_545 (
  .O(mux_o_545),
  .I0(mux_o_290),
  .I1(mux_o_291),
  .S0(ad[5])
);
MUX2 mux_inst_546 (
  .O(mux_o_546),
  .I0(mux_o_292),
  .I1(mux_o_293),
  .S0(ad[5])
);
MUX2 mux_inst_547 (
  .O(mux_o_547),
  .I0(mux_o_294),
  .I1(mux_o_295),
  .S0(ad[5])
);
MUX2 mux_inst_548 (
  .O(mux_o_548),
  .I0(mux_o_296),
  .I1(mux_o_297),
  .S0(ad[5])
);
MUX2 mux_inst_549 (
  .O(mux_o_549),
  .I0(mux_o_298),
  .I1(mux_o_299),
  .S0(ad[5])
);
MUX2 mux_inst_550 (
  .O(mux_o_550),
  .I0(mux_o_300),
  .I1(mux_o_301),
  .S0(ad[5])
);
MUX2 mux_inst_551 (
  .O(mux_o_551),
  .I0(mux_o_302),
  .I1(mux_o_303),
  .S0(ad[5])
);
MUX2 mux_inst_552 (
  .O(mux_o_552),
  .I0(mux_o_304),
  .I1(mux_o_305),
  .S0(ad[5])
);
MUX2 mux_inst_553 (
  .O(mux_o_553),
  .I0(mux_o_306),
  .I1(mux_o_307),
  .S0(ad[5])
);
MUX2 mux_inst_554 (
  .O(mux_o_554),
  .I0(mux_o_308),
  .I1(mux_o_309),
  .S0(ad[5])
);
MUX2 mux_inst_555 (
  .O(mux_o_555),
  .I0(mux_o_310),
  .I1(mux_o_311),
  .S0(ad[5])
);
MUX2 mux_inst_556 (
  .O(mux_o_556),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(ad[5])
);
MUX2 mux_inst_557 (
  .O(mux_o_557),
  .I0(mux_o_314),
  .I1(mux_o_315),
  .S0(ad[5])
);
MUX2 mux_inst_558 (
  .O(mux_o_558),
  .I0(mux_o_316),
  .I1(mux_o_317),
  .S0(ad[5])
);
MUX2 mux_inst_559 (
  .O(mux_o_559),
  .I0(mux_o_318),
  .I1(mux_o_319),
  .S0(ad[5])
);
MUX2 mux_inst_560 (
  .O(mux_o_560),
  .I0(mux_o_320),
  .I1(mux_o_321),
  .S0(ad[5])
);
MUX2 mux_inst_561 (
  .O(mux_o_561),
  .I0(mux_o_322),
  .I1(mux_o_323),
  .S0(ad[5])
);
MUX2 mux_inst_562 (
  .O(mux_o_562),
  .I0(mux_o_324),
  .I1(mux_o_325),
  .S0(ad[5])
);
MUX2 mux_inst_563 (
  .O(mux_o_563),
  .I0(mux_o_326),
  .I1(mux_o_327),
  .S0(ad[5])
);
MUX2 mux_inst_564 (
  .O(mux_o_564),
  .I0(mux_o_328),
  .I1(mux_o_329),
  .S0(ad[5])
);
MUX2 mux_inst_565 (
  .O(mux_o_565),
  .I0(mux_o_330),
  .I1(mux_o_331),
  .S0(ad[5])
);
MUX2 mux_inst_566 (
  .O(mux_o_566),
  .I0(mux_o_332),
  .I1(mux_o_333),
  .S0(ad[5])
);
MUX2 mux_inst_567 (
  .O(mux_o_567),
  .I0(mux_o_334),
  .I1(mux_o_335),
  .S0(ad[5])
);
MUX2 mux_inst_568 (
  .O(mux_o_568),
  .I0(mux_o_336),
  .I1(mux_o_337),
  .S0(ad[5])
);
MUX2 mux_inst_569 (
  .O(mux_o_569),
  .I0(mux_o_338),
  .I1(mux_o_339),
  .S0(ad[5])
);
MUX2 mux_inst_570 (
  .O(mux_o_570),
  .I0(mux_o_340),
  .I1(mux_o_341),
  .S0(ad[5])
);
MUX2 mux_inst_571 (
  .O(mux_o_571),
  .I0(mux_o_342),
  .I1(mux_o_343),
  .S0(ad[5])
);
MUX2 mux_inst_572 (
  .O(mux_o_572),
  .I0(mux_o_344),
  .I1(mux_o_345),
  .S0(ad[5])
);
MUX2 mux_inst_573 (
  .O(mux_o_573),
  .I0(mux_o_346),
  .I1(mux_o_347),
  .S0(ad[5])
);
MUX2 mux_inst_574 (
  .O(mux_o_574),
  .I0(mux_o_348),
  .I1(mux_o_349),
  .S0(ad[5])
);
MUX2 mux_inst_575 (
  .O(mux_o_575),
  .I0(mux_o_350),
  .I1(mux_o_351),
  .S0(ad[5])
);
MUX2 mux_inst_576 (
  .O(mux_o_576),
  .I0(mux_o_352),
  .I1(mux_o_353),
  .S0(ad[5])
);
MUX2 mux_inst_577 (
  .O(mux_o_577),
  .I0(mux_o_354),
  .I1(mux_o_355),
  .S0(ad[5])
);
MUX2 mux_inst_578 (
  .O(mux_o_578),
  .I0(mux_o_356),
  .I1(mux_o_357),
  .S0(ad[5])
);
MUX2 mux_inst_579 (
  .O(mux_o_579),
  .I0(mux_o_358),
  .I1(mux_o_359),
  .S0(ad[5])
);
MUX2 mux_inst_580 (
  .O(mux_o_580),
  .I0(mux_o_360),
  .I1(mux_o_361),
  .S0(ad[5])
);
MUX2 mux_inst_581 (
  .O(mux_o_581),
  .I0(mux_o_362),
  .I1(mux_o_363),
  .S0(ad[5])
);
MUX2 mux_inst_582 (
  .O(mux_o_582),
  .I0(mux_o_364),
  .I1(mux_o_365),
  .S0(ad[5])
);
MUX2 mux_inst_583 (
  .O(mux_o_583),
  .I0(mux_o_366),
  .I1(mux_o_367),
  .S0(ad[5])
);
MUX2 mux_inst_584 (
  .O(mux_o_584),
  .I0(mux_o_368),
  .I1(mux_o_369),
  .S0(ad[5])
);
MUX2 mux_inst_585 (
  .O(mux_o_585),
  .I0(mux_o_370),
  .I1(mux_o_371),
  .S0(ad[5])
);
MUX2 mux_inst_586 (
  .O(mux_o_586),
  .I0(mux_o_372),
  .I1(mux_o_373),
  .S0(ad[5])
);
MUX2 mux_inst_587 (
  .O(mux_o_587),
  .I0(mux_o_374),
  .I1(mux_o_375),
  .S0(ad[5])
);
MUX2 mux_inst_588 (
  .O(mux_o_588),
  .I0(mux_o_376),
  .I1(mux_o_377),
  .S0(ad[5])
);
MUX2 mux_inst_589 (
  .O(mux_o_589),
  .I0(mux_o_378),
  .I1(mux_o_379),
  .S0(ad[5])
);
MUX2 mux_inst_590 (
  .O(mux_o_590),
  .I0(mux_o_380),
  .I1(mux_o_381),
  .S0(ad[5])
);
MUX2 mux_inst_591 (
  .O(mux_o_591),
  .I0(mux_o_382),
  .I1(mux_o_383),
  .S0(ad[5])
);
MUX2 mux_inst_592 (
  .O(mux_o_592),
  .I0(mux_o_384),
  .I1(mux_o_385),
  .S0(ad[5])
);
MUX2 mux_inst_593 (
  .O(mux_o_593),
  .I0(mux_o_386),
  .I1(mux_o_387),
  .S0(ad[5])
);
MUX2 mux_inst_594 (
  .O(mux_o_594),
  .I0(mux_o_388),
  .I1(mux_o_389),
  .S0(ad[5])
);
MUX2 mux_inst_595 (
  .O(mux_o_595),
  .I0(mux_o_390),
  .I1(mux_o_391),
  .S0(ad[5])
);
MUX2 mux_inst_596 (
  .O(mux_o_596),
  .I0(mux_o_392),
  .I1(mux_o_393),
  .S0(ad[5])
);
MUX2 mux_inst_597 (
  .O(mux_o_597),
  .I0(mux_o_394),
  .I1(mux_o_395),
  .S0(ad[5])
);
MUX2 mux_inst_598 (
  .O(mux_o_598),
  .I0(mux_o_396),
  .I1(mux_o_397),
  .S0(ad[5])
);
MUX2 mux_inst_599 (
  .O(mux_o_599),
  .I0(mux_o_398),
  .I1(mux_o_399),
  .S0(ad[5])
);
MUX2 mux_inst_600 (
  .O(mux_o_600),
  .I0(mux_o_400),
  .I1(mux_o_401),
  .S0(ad[6])
);
MUX2 mux_inst_601 (
  .O(mux_o_601),
  .I0(mux_o_402),
  .I1(mux_o_403),
  .S0(ad[6])
);
MUX2 mux_inst_602 (
  .O(mux_o_602),
  .I0(mux_o_404),
  .I1(mux_o_405),
  .S0(ad[6])
);
MUX2 mux_inst_603 (
  .O(mux_o_603),
  .I0(mux_o_406),
  .I1(mux_o_407),
  .S0(ad[6])
);
MUX2 mux_inst_604 (
  .O(mux_o_604),
  .I0(mux_o_408),
  .I1(mux_o_409),
  .S0(ad[6])
);
MUX2 mux_inst_605 (
  .O(mux_o_605),
  .I0(mux_o_410),
  .I1(mux_o_411),
  .S0(ad[6])
);
MUX2 mux_inst_606 (
  .O(mux_o_606),
  .I0(mux_o_412),
  .I1(mux_o_413),
  .S0(ad[6])
);
MUX2 mux_inst_607 (
  .O(mux_o_607),
  .I0(mux_o_414),
  .I1(mux_o_415),
  .S0(ad[6])
);
MUX2 mux_inst_608 (
  .O(mux_o_608),
  .I0(mux_o_416),
  .I1(mux_o_417),
  .S0(ad[6])
);
MUX2 mux_inst_609 (
  .O(mux_o_609),
  .I0(mux_o_418),
  .I1(mux_o_419),
  .S0(ad[6])
);
MUX2 mux_inst_610 (
  .O(mux_o_610),
  .I0(mux_o_420),
  .I1(mux_o_421),
  .S0(ad[6])
);
MUX2 mux_inst_611 (
  .O(mux_o_611),
  .I0(mux_o_422),
  .I1(mux_o_423),
  .S0(ad[6])
);
MUX2 mux_inst_612 (
  .O(mux_o_612),
  .I0(mux_o_424),
  .I1(mux_o_425),
  .S0(ad[6])
);
MUX2 mux_inst_613 (
  .O(mux_o_613),
  .I0(mux_o_426),
  .I1(mux_o_427),
  .S0(ad[6])
);
MUX2 mux_inst_614 (
  .O(mux_o_614),
  .I0(mux_o_428),
  .I1(mux_o_429),
  .S0(ad[6])
);
MUX2 mux_inst_615 (
  .O(mux_o_615),
  .I0(mux_o_430),
  .I1(mux_o_431),
  .S0(ad[6])
);
MUX2 mux_inst_616 (
  .O(mux_o_616),
  .I0(mux_o_432),
  .I1(mux_o_433),
  .S0(ad[6])
);
MUX2 mux_inst_617 (
  .O(mux_o_617),
  .I0(mux_o_434),
  .I1(mux_o_435),
  .S0(ad[6])
);
MUX2 mux_inst_618 (
  .O(mux_o_618),
  .I0(mux_o_436),
  .I1(mux_o_437),
  .S0(ad[6])
);
MUX2 mux_inst_619 (
  .O(mux_o_619),
  .I0(mux_o_438),
  .I1(mux_o_439),
  .S0(ad[6])
);
MUX2 mux_inst_620 (
  .O(mux_o_620),
  .I0(mux_o_440),
  .I1(mux_o_441),
  .S0(ad[6])
);
MUX2 mux_inst_621 (
  .O(mux_o_621),
  .I0(mux_o_442),
  .I1(mux_o_443),
  .S0(ad[6])
);
MUX2 mux_inst_622 (
  .O(mux_o_622),
  .I0(mux_o_444),
  .I1(mux_o_445),
  .S0(ad[6])
);
MUX2 mux_inst_623 (
  .O(mux_o_623),
  .I0(mux_o_446),
  .I1(mux_o_447),
  .S0(ad[6])
);
MUX2 mux_inst_624 (
  .O(mux_o_624),
  .I0(mux_o_448),
  .I1(mux_o_449),
  .S0(ad[6])
);
MUX2 mux_inst_625 (
  .O(mux_o_625),
  .I0(mux_o_450),
  .I1(mux_o_451),
  .S0(ad[6])
);
MUX2 mux_inst_626 (
  .O(mux_o_626),
  .I0(mux_o_452),
  .I1(mux_o_453),
  .S0(ad[6])
);
MUX2 mux_inst_627 (
  .O(mux_o_627),
  .I0(mux_o_454),
  .I1(mux_o_455),
  .S0(ad[6])
);
MUX2 mux_inst_628 (
  .O(mux_o_628),
  .I0(mux_o_456),
  .I1(mux_o_457),
  .S0(ad[6])
);
MUX2 mux_inst_629 (
  .O(mux_o_629),
  .I0(mux_o_458),
  .I1(mux_o_459),
  .S0(ad[6])
);
MUX2 mux_inst_630 (
  .O(mux_o_630),
  .I0(mux_o_460),
  .I1(mux_o_461),
  .S0(ad[6])
);
MUX2 mux_inst_631 (
  .O(mux_o_631),
  .I0(mux_o_462),
  .I1(mux_o_463),
  .S0(ad[6])
);
MUX2 mux_inst_632 (
  .O(mux_o_632),
  .I0(mux_o_464),
  .I1(mux_o_465),
  .S0(ad[6])
);
MUX2 mux_inst_633 (
  .O(mux_o_633),
  .I0(mux_o_466),
  .I1(mux_o_467),
  .S0(ad[6])
);
MUX2 mux_inst_634 (
  .O(mux_o_634),
  .I0(mux_o_468),
  .I1(mux_o_469),
  .S0(ad[6])
);
MUX2 mux_inst_635 (
  .O(mux_o_635),
  .I0(mux_o_470),
  .I1(mux_o_471),
  .S0(ad[6])
);
MUX2 mux_inst_636 (
  .O(mux_o_636),
  .I0(mux_o_472),
  .I1(mux_o_473),
  .S0(ad[6])
);
MUX2 mux_inst_637 (
  .O(mux_o_637),
  .I0(mux_o_474),
  .I1(mux_o_475),
  .S0(ad[6])
);
MUX2 mux_inst_638 (
  .O(mux_o_638),
  .I0(mux_o_476),
  .I1(mux_o_477),
  .S0(ad[6])
);
MUX2 mux_inst_639 (
  .O(mux_o_639),
  .I0(mux_o_478),
  .I1(mux_o_479),
  .S0(ad[6])
);
MUX2 mux_inst_640 (
  .O(mux_o_640),
  .I0(mux_o_480),
  .I1(mux_o_481),
  .S0(ad[6])
);
MUX2 mux_inst_641 (
  .O(mux_o_641),
  .I0(mux_o_482),
  .I1(mux_o_483),
  .S0(ad[6])
);
MUX2 mux_inst_642 (
  .O(mux_o_642),
  .I0(mux_o_484),
  .I1(mux_o_485),
  .S0(ad[6])
);
MUX2 mux_inst_643 (
  .O(mux_o_643),
  .I0(mux_o_486),
  .I1(mux_o_487),
  .S0(ad[6])
);
MUX2 mux_inst_644 (
  .O(mux_o_644),
  .I0(mux_o_488),
  .I1(mux_o_489),
  .S0(ad[6])
);
MUX2 mux_inst_645 (
  .O(mux_o_645),
  .I0(mux_o_490),
  .I1(mux_o_491),
  .S0(ad[6])
);
MUX2 mux_inst_646 (
  .O(mux_o_646),
  .I0(mux_o_492),
  .I1(mux_o_493),
  .S0(ad[6])
);
MUX2 mux_inst_647 (
  .O(mux_o_647),
  .I0(mux_o_494),
  .I1(mux_o_495),
  .S0(ad[6])
);
MUX2 mux_inst_648 (
  .O(mux_o_648),
  .I0(mux_o_496),
  .I1(mux_o_497),
  .S0(ad[6])
);
MUX2 mux_inst_649 (
  .O(mux_o_649),
  .I0(mux_o_498),
  .I1(mux_o_499),
  .S0(ad[6])
);
MUX2 mux_inst_650 (
  .O(mux_o_650),
  .I0(mux_o_500),
  .I1(mux_o_501),
  .S0(ad[6])
);
MUX2 mux_inst_651 (
  .O(mux_o_651),
  .I0(mux_o_502),
  .I1(mux_o_503),
  .S0(ad[6])
);
MUX2 mux_inst_652 (
  .O(mux_o_652),
  .I0(mux_o_504),
  .I1(mux_o_505),
  .S0(ad[6])
);
MUX2 mux_inst_653 (
  .O(mux_o_653),
  .I0(mux_o_506),
  .I1(mux_o_507),
  .S0(ad[6])
);
MUX2 mux_inst_654 (
  .O(mux_o_654),
  .I0(mux_o_508),
  .I1(mux_o_509),
  .S0(ad[6])
);
MUX2 mux_inst_655 (
  .O(mux_o_655),
  .I0(mux_o_510),
  .I1(mux_o_511),
  .S0(ad[6])
);
MUX2 mux_inst_656 (
  .O(mux_o_656),
  .I0(mux_o_512),
  .I1(mux_o_513),
  .S0(ad[6])
);
MUX2 mux_inst_657 (
  .O(mux_o_657),
  .I0(mux_o_514),
  .I1(mux_o_515),
  .S0(ad[6])
);
MUX2 mux_inst_658 (
  .O(mux_o_658),
  .I0(mux_o_516),
  .I1(mux_o_517),
  .S0(ad[6])
);
MUX2 mux_inst_659 (
  .O(mux_o_659),
  .I0(mux_o_518),
  .I1(mux_o_519),
  .S0(ad[6])
);
MUX2 mux_inst_660 (
  .O(mux_o_660),
  .I0(mux_o_520),
  .I1(mux_o_521),
  .S0(ad[6])
);
MUX2 mux_inst_661 (
  .O(mux_o_661),
  .I0(mux_o_522),
  .I1(mux_o_523),
  .S0(ad[6])
);
MUX2 mux_inst_662 (
  .O(mux_o_662),
  .I0(mux_o_524),
  .I1(mux_o_525),
  .S0(ad[6])
);
MUX2 mux_inst_663 (
  .O(mux_o_663),
  .I0(mux_o_526),
  .I1(mux_o_527),
  .S0(ad[6])
);
MUX2 mux_inst_664 (
  .O(mux_o_664),
  .I0(mux_o_528),
  .I1(mux_o_529),
  .S0(ad[6])
);
MUX2 mux_inst_665 (
  .O(mux_o_665),
  .I0(mux_o_530),
  .I1(mux_o_531),
  .S0(ad[6])
);
MUX2 mux_inst_666 (
  .O(mux_o_666),
  .I0(mux_o_532),
  .I1(mux_o_533),
  .S0(ad[6])
);
MUX2 mux_inst_667 (
  .O(mux_o_667),
  .I0(mux_o_534),
  .I1(mux_o_535),
  .S0(ad[6])
);
MUX2 mux_inst_668 (
  .O(mux_o_668),
  .I0(mux_o_536),
  .I1(mux_o_537),
  .S0(ad[6])
);
MUX2 mux_inst_669 (
  .O(mux_o_669),
  .I0(mux_o_538),
  .I1(mux_o_539),
  .S0(ad[6])
);
MUX2 mux_inst_670 (
  .O(mux_o_670),
  .I0(mux_o_540),
  .I1(mux_o_541),
  .S0(ad[6])
);
MUX2 mux_inst_671 (
  .O(mux_o_671),
  .I0(mux_o_542),
  .I1(mux_o_543),
  .S0(ad[6])
);
MUX2 mux_inst_672 (
  .O(mux_o_672),
  .I0(mux_o_544),
  .I1(mux_o_545),
  .S0(ad[6])
);
MUX2 mux_inst_673 (
  .O(mux_o_673),
  .I0(mux_o_546),
  .I1(mux_o_547),
  .S0(ad[6])
);
MUX2 mux_inst_674 (
  .O(mux_o_674),
  .I0(mux_o_548),
  .I1(mux_o_549),
  .S0(ad[6])
);
MUX2 mux_inst_675 (
  .O(mux_o_675),
  .I0(mux_o_550),
  .I1(mux_o_551),
  .S0(ad[6])
);
MUX2 mux_inst_676 (
  .O(mux_o_676),
  .I0(mux_o_552),
  .I1(mux_o_553),
  .S0(ad[6])
);
MUX2 mux_inst_677 (
  .O(mux_o_677),
  .I0(mux_o_554),
  .I1(mux_o_555),
  .S0(ad[6])
);
MUX2 mux_inst_678 (
  .O(mux_o_678),
  .I0(mux_o_556),
  .I1(mux_o_557),
  .S0(ad[6])
);
MUX2 mux_inst_679 (
  .O(mux_o_679),
  .I0(mux_o_558),
  .I1(mux_o_559),
  .S0(ad[6])
);
MUX2 mux_inst_680 (
  .O(mux_o_680),
  .I0(mux_o_560),
  .I1(mux_o_561),
  .S0(ad[6])
);
MUX2 mux_inst_681 (
  .O(mux_o_681),
  .I0(mux_o_562),
  .I1(mux_o_563),
  .S0(ad[6])
);
MUX2 mux_inst_682 (
  .O(mux_o_682),
  .I0(mux_o_564),
  .I1(mux_o_565),
  .S0(ad[6])
);
MUX2 mux_inst_683 (
  .O(mux_o_683),
  .I0(mux_o_566),
  .I1(mux_o_567),
  .S0(ad[6])
);
MUX2 mux_inst_684 (
  .O(mux_o_684),
  .I0(mux_o_568),
  .I1(mux_o_569),
  .S0(ad[6])
);
MUX2 mux_inst_685 (
  .O(mux_o_685),
  .I0(mux_o_570),
  .I1(mux_o_571),
  .S0(ad[6])
);
MUX2 mux_inst_686 (
  .O(mux_o_686),
  .I0(mux_o_572),
  .I1(mux_o_573),
  .S0(ad[6])
);
MUX2 mux_inst_687 (
  .O(mux_o_687),
  .I0(mux_o_574),
  .I1(mux_o_575),
  .S0(ad[6])
);
MUX2 mux_inst_688 (
  .O(mux_o_688),
  .I0(mux_o_576),
  .I1(mux_o_577),
  .S0(ad[6])
);
MUX2 mux_inst_689 (
  .O(mux_o_689),
  .I0(mux_o_578),
  .I1(mux_o_579),
  .S0(ad[6])
);
MUX2 mux_inst_690 (
  .O(mux_o_690),
  .I0(mux_o_580),
  .I1(mux_o_581),
  .S0(ad[6])
);
MUX2 mux_inst_691 (
  .O(mux_o_691),
  .I0(mux_o_582),
  .I1(mux_o_583),
  .S0(ad[6])
);
MUX2 mux_inst_692 (
  .O(mux_o_692),
  .I0(mux_o_584),
  .I1(mux_o_585),
  .S0(ad[6])
);
MUX2 mux_inst_693 (
  .O(mux_o_693),
  .I0(mux_o_586),
  .I1(mux_o_587),
  .S0(ad[6])
);
MUX2 mux_inst_694 (
  .O(mux_o_694),
  .I0(mux_o_588),
  .I1(mux_o_589),
  .S0(ad[6])
);
MUX2 mux_inst_695 (
  .O(mux_o_695),
  .I0(mux_o_590),
  .I1(mux_o_591),
  .S0(ad[6])
);
MUX2 mux_inst_696 (
  .O(mux_o_696),
  .I0(mux_o_592),
  .I1(mux_o_593),
  .S0(ad[6])
);
MUX2 mux_inst_697 (
  .O(mux_o_697),
  .I0(mux_o_594),
  .I1(mux_o_595),
  .S0(ad[6])
);
MUX2 mux_inst_698 (
  .O(mux_o_698),
  .I0(mux_o_596),
  .I1(mux_o_597),
  .S0(ad[6])
);
MUX2 mux_inst_699 (
  .O(mux_o_699),
  .I0(mux_o_598),
  .I1(mux_o_599),
  .S0(ad[6])
);
MUX2 mux_inst_700 (
  .O(mux_o_700),
  .I0(mux_o_600),
  .I1(mux_o_601),
  .S0(ad[7])
);
MUX2 mux_inst_701 (
  .O(mux_o_701),
  .I0(mux_o_602),
  .I1(mux_o_603),
  .S0(ad[7])
);
MUX2 mux_inst_702 (
  .O(mux_o_702),
  .I0(mux_o_604),
  .I1(mux_o_605),
  .S0(ad[7])
);
MUX2 mux_inst_703 (
  .O(mux_o_703),
  .I0(mux_o_606),
  .I1(mux_o_607),
  .S0(ad[7])
);
MUX2 mux_inst_704 (
  .O(mux_o_704),
  .I0(mux_o_608),
  .I1(mux_o_609),
  .S0(ad[7])
);
MUX2 mux_inst_705 (
  .O(mux_o_705),
  .I0(mux_o_610),
  .I1(mux_o_611),
  .S0(ad[7])
);
MUX2 mux_inst_706 (
  .O(mux_o_706),
  .I0(mux_o_612),
  .I1(mux_o_613),
  .S0(ad[7])
);
MUX2 mux_inst_707 (
  .O(mux_o_707),
  .I0(mux_o_614),
  .I1(mux_o_615),
  .S0(ad[7])
);
MUX2 mux_inst_708 (
  .O(mux_o_708),
  .I0(mux_o_616),
  .I1(mux_o_617),
  .S0(ad[7])
);
MUX2 mux_inst_709 (
  .O(mux_o_709),
  .I0(mux_o_618),
  .I1(mux_o_619),
  .S0(ad[7])
);
MUX2 mux_inst_710 (
  .O(mux_o_710),
  .I0(mux_o_620),
  .I1(mux_o_621),
  .S0(ad[7])
);
MUX2 mux_inst_711 (
  .O(mux_o_711),
  .I0(mux_o_622),
  .I1(mux_o_623),
  .S0(ad[7])
);
MUX2 mux_inst_712 (
  .O(mux_o_712),
  .I0(mux_o_624),
  .I1(mux_o_625),
  .S0(ad[7])
);
MUX2 mux_inst_713 (
  .O(mux_o_713),
  .I0(mux_o_626),
  .I1(mux_o_627),
  .S0(ad[7])
);
MUX2 mux_inst_714 (
  .O(mux_o_714),
  .I0(mux_o_628),
  .I1(mux_o_629),
  .S0(ad[7])
);
MUX2 mux_inst_715 (
  .O(mux_o_715),
  .I0(mux_o_630),
  .I1(mux_o_631),
  .S0(ad[7])
);
MUX2 mux_inst_716 (
  .O(mux_o_716),
  .I0(mux_o_632),
  .I1(mux_o_633),
  .S0(ad[7])
);
MUX2 mux_inst_717 (
  .O(mux_o_717),
  .I0(mux_o_634),
  .I1(mux_o_635),
  .S0(ad[7])
);
MUX2 mux_inst_718 (
  .O(mux_o_718),
  .I0(mux_o_636),
  .I1(mux_o_637),
  .S0(ad[7])
);
MUX2 mux_inst_719 (
  .O(mux_o_719),
  .I0(mux_o_638),
  .I1(mux_o_639),
  .S0(ad[7])
);
MUX2 mux_inst_720 (
  .O(mux_o_720),
  .I0(mux_o_640),
  .I1(mux_o_641),
  .S0(ad[7])
);
MUX2 mux_inst_721 (
  .O(mux_o_721),
  .I0(mux_o_642),
  .I1(mux_o_643),
  .S0(ad[7])
);
MUX2 mux_inst_722 (
  .O(mux_o_722),
  .I0(mux_o_644),
  .I1(mux_o_645),
  .S0(ad[7])
);
MUX2 mux_inst_723 (
  .O(mux_o_723),
  .I0(mux_o_646),
  .I1(mux_o_647),
  .S0(ad[7])
);
MUX2 mux_inst_724 (
  .O(mux_o_724),
  .I0(mux_o_648),
  .I1(mux_o_649),
  .S0(ad[7])
);
MUX2 mux_inst_725 (
  .O(mux_o_725),
  .I0(mux_o_650),
  .I1(mux_o_651),
  .S0(ad[7])
);
MUX2 mux_inst_726 (
  .O(mux_o_726),
  .I0(mux_o_652),
  .I1(mux_o_653),
  .S0(ad[7])
);
MUX2 mux_inst_727 (
  .O(mux_o_727),
  .I0(mux_o_654),
  .I1(mux_o_655),
  .S0(ad[7])
);
MUX2 mux_inst_728 (
  .O(mux_o_728),
  .I0(mux_o_656),
  .I1(mux_o_657),
  .S0(ad[7])
);
MUX2 mux_inst_729 (
  .O(mux_o_729),
  .I0(mux_o_658),
  .I1(mux_o_659),
  .S0(ad[7])
);
MUX2 mux_inst_730 (
  .O(mux_o_730),
  .I0(mux_o_660),
  .I1(mux_o_661),
  .S0(ad[7])
);
MUX2 mux_inst_731 (
  .O(mux_o_731),
  .I0(mux_o_662),
  .I1(mux_o_663),
  .S0(ad[7])
);
MUX2 mux_inst_732 (
  .O(mux_o_732),
  .I0(mux_o_664),
  .I1(mux_o_665),
  .S0(ad[7])
);
MUX2 mux_inst_733 (
  .O(mux_o_733),
  .I0(mux_o_666),
  .I1(mux_o_667),
  .S0(ad[7])
);
MUX2 mux_inst_734 (
  .O(mux_o_734),
  .I0(mux_o_668),
  .I1(mux_o_669),
  .S0(ad[7])
);
MUX2 mux_inst_735 (
  .O(mux_o_735),
  .I0(mux_o_670),
  .I1(mux_o_671),
  .S0(ad[7])
);
MUX2 mux_inst_736 (
  .O(mux_o_736),
  .I0(mux_o_672),
  .I1(mux_o_673),
  .S0(ad[7])
);
MUX2 mux_inst_737 (
  .O(mux_o_737),
  .I0(mux_o_674),
  .I1(mux_o_675),
  .S0(ad[7])
);
MUX2 mux_inst_738 (
  .O(mux_o_738),
  .I0(mux_o_676),
  .I1(mux_o_677),
  .S0(ad[7])
);
MUX2 mux_inst_739 (
  .O(mux_o_739),
  .I0(mux_o_678),
  .I1(mux_o_679),
  .S0(ad[7])
);
MUX2 mux_inst_740 (
  .O(mux_o_740),
  .I0(mux_o_680),
  .I1(mux_o_681),
  .S0(ad[7])
);
MUX2 mux_inst_741 (
  .O(mux_o_741),
  .I0(mux_o_682),
  .I1(mux_o_683),
  .S0(ad[7])
);
MUX2 mux_inst_742 (
  .O(mux_o_742),
  .I0(mux_o_684),
  .I1(mux_o_685),
  .S0(ad[7])
);
MUX2 mux_inst_743 (
  .O(mux_o_743),
  .I0(mux_o_686),
  .I1(mux_o_687),
  .S0(ad[7])
);
MUX2 mux_inst_744 (
  .O(mux_o_744),
  .I0(mux_o_688),
  .I1(mux_o_689),
  .S0(ad[7])
);
MUX2 mux_inst_745 (
  .O(mux_o_745),
  .I0(mux_o_690),
  .I1(mux_o_691),
  .S0(ad[7])
);
MUX2 mux_inst_746 (
  .O(mux_o_746),
  .I0(mux_o_692),
  .I1(mux_o_693),
  .S0(ad[7])
);
MUX2 mux_inst_747 (
  .O(mux_o_747),
  .I0(mux_o_694),
  .I1(mux_o_695),
  .S0(ad[7])
);
MUX2 mux_inst_748 (
  .O(mux_o_748),
  .I0(mux_o_696),
  .I1(mux_o_697),
  .S0(ad[7])
);
MUX2 mux_inst_749 (
  .O(mux_o_749),
  .I0(mux_o_698),
  .I1(mux_o_699),
  .S0(ad[7])
);
MUX2 mux_inst_750 (
  .O(mux_o_750),
  .I0(mux_o_700),
  .I1(mux_o_701),
  .S0(ad[8])
);
MUX2 mux_inst_751 (
  .O(mux_o_751),
  .I0(mux_o_702),
  .I1(mux_o_703),
  .S0(ad[8])
);
MUX2 mux_inst_752 (
  .O(mux_o_752),
  .I0(mux_o_704),
  .I1(mux_o_705),
  .S0(ad[8])
);
MUX2 mux_inst_753 (
  .O(mux_o_753),
  .I0(mux_o_706),
  .I1(mux_o_707),
  .S0(ad[8])
);
MUX2 mux_inst_754 (
  .O(mux_o_754),
  .I0(mux_o_708),
  .I1(mux_o_709),
  .S0(ad[8])
);
MUX2 mux_inst_755 (
  .O(mux_o_755),
  .I0(mux_o_710),
  .I1(mux_o_711),
  .S0(ad[8])
);
MUX2 mux_inst_756 (
  .O(mux_o_756),
  .I0(mux_o_712),
  .I1(mux_o_713),
  .S0(ad[8])
);
MUX2 mux_inst_757 (
  .O(mux_o_757),
  .I0(mux_o_714),
  .I1(mux_o_715),
  .S0(ad[8])
);
MUX2 mux_inst_758 (
  .O(mux_o_758),
  .I0(mux_o_716),
  .I1(mux_o_717),
  .S0(ad[8])
);
MUX2 mux_inst_759 (
  .O(mux_o_759),
  .I0(mux_o_718),
  .I1(mux_o_719),
  .S0(ad[8])
);
MUX2 mux_inst_760 (
  .O(mux_o_760),
  .I0(mux_o_720),
  .I1(mux_o_721),
  .S0(ad[8])
);
MUX2 mux_inst_761 (
  .O(mux_o_761),
  .I0(mux_o_722),
  .I1(mux_o_723),
  .S0(ad[8])
);
MUX2 mux_inst_762 (
  .O(mux_o_762),
  .I0(mux_o_724),
  .I1(mux_o_725),
  .S0(ad[8])
);
MUX2 mux_inst_763 (
  .O(mux_o_763),
  .I0(mux_o_726),
  .I1(mux_o_727),
  .S0(ad[8])
);
MUX2 mux_inst_764 (
  .O(mux_o_764),
  .I0(mux_o_728),
  .I1(mux_o_729),
  .S0(ad[8])
);
MUX2 mux_inst_765 (
  .O(mux_o_765),
  .I0(mux_o_730),
  .I1(mux_o_731),
  .S0(ad[8])
);
MUX2 mux_inst_766 (
  .O(mux_o_766),
  .I0(mux_o_732),
  .I1(mux_o_733),
  .S0(ad[8])
);
MUX2 mux_inst_767 (
  .O(mux_o_767),
  .I0(mux_o_734),
  .I1(mux_o_735),
  .S0(ad[8])
);
MUX2 mux_inst_768 (
  .O(mux_o_768),
  .I0(mux_o_736),
  .I1(mux_o_737),
  .S0(ad[8])
);
MUX2 mux_inst_769 (
  .O(mux_o_769),
  .I0(mux_o_738),
  .I1(mux_o_739),
  .S0(ad[8])
);
MUX2 mux_inst_770 (
  .O(mux_o_770),
  .I0(mux_o_740),
  .I1(mux_o_741),
  .S0(ad[8])
);
MUX2 mux_inst_771 (
  .O(mux_o_771),
  .I0(mux_o_742),
  .I1(mux_o_743),
  .S0(ad[8])
);
MUX2 mux_inst_772 (
  .O(mux_o_772),
  .I0(mux_o_744),
  .I1(mux_o_745),
  .S0(ad[8])
);
MUX2 mux_inst_773 (
  .O(mux_o_773),
  .I0(mux_o_746),
  .I1(mux_o_747),
  .S0(ad[8])
);
MUX2 mux_inst_774 (
  .O(mux_o_774),
  .I0(mux_o_748),
  .I1(mux_o_749),
  .S0(ad[8])
);
MUX2 mux_inst_775 (
  .O(mux_o_775),
  .I0(mux_o_750),
  .I1(mux_o_751),
  .S0(ad[9])
);
MUX2 mux_inst_776 (
  .O(mux_o_776),
  .I0(mux_o_752),
  .I1(mux_o_753),
  .S0(ad[9])
);
MUX2 mux_inst_777 (
  .O(mux_o_777),
  .I0(mux_o_754),
  .I1(mux_o_755),
  .S0(ad[9])
);
MUX2 mux_inst_778 (
  .O(mux_o_778),
  .I0(mux_o_756),
  .I1(mux_o_757),
  .S0(ad[9])
);
MUX2 mux_inst_779 (
  .O(mux_o_779),
  .I0(mux_o_758),
  .I1(mux_o_759),
  .S0(ad[9])
);
MUX2 mux_inst_780 (
  .O(mux_o_780),
  .I0(mux_o_760),
  .I1(mux_o_761),
  .S0(ad[9])
);
MUX2 mux_inst_781 (
  .O(mux_o_781),
  .I0(mux_o_762),
  .I1(mux_o_763),
  .S0(ad[9])
);
MUX2 mux_inst_782 (
  .O(mux_o_782),
  .I0(mux_o_764),
  .I1(mux_o_765),
  .S0(ad[9])
);
MUX2 mux_inst_783 (
  .O(mux_o_783),
  .I0(mux_o_766),
  .I1(mux_o_767),
  .S0(ad[9])
);
MUX2 mux_inst_784 (
  .O(mux_o_784),
  .I0(mux_o_768),
  .I1(mux_o_769),
  .S0(ad[9])
);
MUX2 mux_inst_785 (
  .O(mux_o_785),
  .I0(mux_o_770),
  .I1(mux_o_771),
  .S0(ad[9])
);
MUX2 mux_inst_786 (
  .O(mux_o_786),
  .I0(mux_o_772),
  .I1(mux_o_773),
  .S0(ad[9])
);
MUX2 mux_inst_788 (
  .O(mux_o_788),
  .I0(mux_o_775),
  .I1(mux_o_776),
  .S0(ad[10])
);
MUX2 mux_inst_789 (
  .O(mux_o_789),
  .I0(mux_o_777),
  .I1(mux_o_778),
  .S0(ad[10])
);
MUX2 mux_inst_790 (
  .O(mux_o_790),
  .I0(mux_o_779),
  .I1(mux_o_780),
  .S0(ad[10])
);
MUX2 mux_inst_791 (
  .O(mux_o_791),
  .I0(mux_o_781),
  .I1(mux_o_782),
  .S0(ad[10])
);
MUX2 mux_inst_792 (
  .O(mux_o_792),
  .I0(mux_o_783),
  .I1(mux_o_784),
  .S0(ad[10])
);
MUX2 mux_inst_793 (
  .O(mux_o_793),
  .I0(mux_o_785),
  .I1(mux_o_786),
  .S0(ad[10])
);
MUX2 mux_inst_795 (
  .O(mux_o_795),
  .I0(mux_o_788),
  .I1(mux_o_789),
  .S0(ad[11])
);
MUX2 mux_inst_796 (
  .O(mux_o_796),
  .I0(mux_o_790),
  .I1(mux_o_791),
  .S0(ad[11])
);
MUX2 mux_inst_797 (
  .O(mux_o_797),
  .I0(mux_o_792),
  .I1(mux_o_793),
  .S0(ad[11])
);
MUX2 mux_inst_799 (
  .O(mux_o_799),
  .I0(mux_o_795),
  .I1(mux_o_796),
  .S0(ad[12])
);
MUX2 mux_inst_800 (
  .O(mux_o_800),
  .I0(mux_o_797),
  .I1(mux_o_774),
  .S0(ad[12])
);
MUX2 mux_inst_801 (
  .O(dout[0]),
  .I0(mux_o_799),
  .I1(mux_o_800),
  .S0(ad[13])
);
MUX2 mux_inst_802 (
  .O(mux_o_802),
  .I0(ram16s_inst_0_dout[1]),
  .I1(ram16s_inst_1_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_803 (
  .O(mux_o_803),
  .I0(ram16s_inst_2_dout[1]),
  .I1(ram16s_inst_3_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_804 (
  .O(mux_o_804),
  .I0(ram16s_inst_4_dout[1]),
  .I1(ram16s_inst_5_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_805 (
  .O(mux_o_805),
  .I0(ram16s_inst_6_dout[1]),
  .I1(ram16s_inst_7_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_806 (
  .O(mux_o_806),
  .I0(ram16s_inst_8_dout[1]),
  .I1(ram16s_inst_9_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_807 (
  .O(mux_o_807),
  .I0(ram16s_inst_10_dout[1]),
  .I1(ram16s_inst_11_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_808 (
  .O(mux_o_808),
  .I0(ram16s_inst_12_dout[1]),
  .I1(ram16s_inst_13_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_809 (
  .O(mux_o_809),
  .I0(ram16s_inst_14_dout[1]),
  .I1(ram16s_inst_15_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_810 (
  .O(mux_o_810),
  .I0(ram16s_inst_16_dout[1]),
  .I1(ram16s_inst_17_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_811 (
  .O(mux_o_811),
  .I0(ram16s_inst_18_dout[1]),
  .I1(ram16s_inst_19_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_812 (
  .O(mux_o_812),
  .I0(ram16s_inst_20_dout[1]),
  .I1(ram16s_inst_21_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_813 (
  .O(mux_o_813),
  .I0(ram16s_inst_22_dout[1]),
  .I1(ram16s_inst_23_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_814 (
  .O(mux_o_814),
  .I0(ram16s_inst_24_dout[1]),
  .I1(ram16s_inst_25_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_815 (
  .O(mux_o_815),
  .I0(ram16s_inst_26_dout[1]),
  .I1(ram16s_inst_27_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_816 (
  .O(mux_o_816),
  .I0(ram16s_inst_28_dout[1]),
  .I1(ram16s_inst_29_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_817 (
  .O(mux_o_817),
  .I0(ram16s_inst_30_dout[1]),
  .I1(ram16s_inst_31_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_818 (
  .O(mux_o_818),
  .I0(ram16s_inst_32_dout[1]),
  .I1(ram16s_inst_33_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_819 (
  .O(mux_o_819),
  .I0(ram16s_inst_34_dout[1]),
  .I1(ram16s_inst_35_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_820 (
  .O(mux_o_820),
  .I0(ram16s_inst_36_dout[1]),
  .I1(ram16s_inst_37_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_821 (
  .O(mux_o_821),
  .I0(ram16s_inst_38_dout[1]),
  .I1(ram16s_inst_39_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_822 (
  .O(mux_o_822),
  .I0(ram16s_inst_40_dout[1]),
  .I1(ram16s_inst_41_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_823 (
  .O(mux_o_823),
  .I0(ram16s_inst_42_dout[1]),
  .I1(ram16s_inst_43_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_824 (
  .O(mux_o_824),
  .I0(ram16s_inst_44_dout[1]),
  .I1(ram16s_inst_45_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_825 (
  .O(mux_o_825),
  .I0(ram16s_inst_46_dout[1]),
  .I1(ram16s_inst_47_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_826 (
  .O(mux_o_826),
  .I0(ram16s_inst_48_dout[1]),
  .I1(ram16s_inst_49_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_827 (
  .O(mux_o_827),
  .I0(ram16s_inst_50_dout[1]),
  .I1(ram16s_inst_51_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_828 (
  .O(mux_o_828),
  .I0(ram16s_inst_52_dout[1]),
  .I1(ram16s_inst_53_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_829 (
  .O(mux_o_829),
  .I0(ram16s_inst_54_dout[1]),
  .I1(ram16s_inst_55_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_830 (
  .O(mux_o_830),
  .I0(ram16s_inst_56_dout[1]),
  .I1(ram16s_inst_57_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_831 (
  .O(mux_o_831),
  .I0(ram16s_inst_58_dout[1]),
  .I1(ram16s_inst_59_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_832 (
  .O(mux_o_832),
  .I0(ram16s_inst_60_dout[1]),
  .I1(ram16s_inst_61_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_833 (
  .O(mux_o_833),
  .I0(ram16s_inst_62_dout[1]),
  .I1(ram16s_inst_63_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_834 (
  .O(mux_o_834),
  .I0(ram16s_inst_64_dout[1]),
  .I1(ram16s_inst_65_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_835 (
  .O(mux_o_835),
  .I0(ram16s_inst_66_dout[1]),
  .I1(ram16s_inst_67_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_836 (
  .O(mux_o_836),
  .I0(ram16s_inst_68_dout[1]),
  .I1(ram16s_inst_69_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_837 (
  .O(mux_o_837),
  .I0(ram16s_inst_70_dout[1]),
  .I1(ram16s_inst_71_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_838 (
  .O(mux_o_838),
  .I0(ram16s_inst_72_dout[1]),
  .I1(ram16s_inst_73_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_839 (
  .O(mux_o_839),
  .I0(ram16s_inst_74_dout[1]),
  .I1(ram16s_inst_75_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_840 (
  .O(mux_o_840),
  .I0(ram16s_inst_76_dout[1]),
  .I1(ram16s_inst_77_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_841 (
  .O(mux_o_841),
  .I0(ram16s_inst_78_dout[1]),
  .I1(ram16s_inst_79_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_842 (
  .O(mux_o_842),
  .I0(ram16s_inst_80_dout[1]),
  .I1(ram16s_inst_81_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_843 (
  .O(mux_o_843),
  .I0(ram16s_inst_82_dout[1]),
  .I1(ram16s_inst_83_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_844 (
  .O(mux_o_844),
  .I0(ram16s_inst_84_dout[1]),
  .I1(ram16s_inst_85_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_845 (
  .O(mux_o_845),
  .I0(ram16s_inst_86_dout[1]),
  .I1(ram16s_inst_87_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_846 (
  .O(mux_o_846),
  .I0(ram16s_inst_88_dout[1]),
  .I1(ram16s_inst_89_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_847 (
  .O(mux_o_847),
  .I0(ram16s_inst_90_dout[1]),
  .I1(ram16s_inst_91_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_848 (
  .O(mux_o_848),
  .I0(ram16s_inst_92_dout[1]),
  .I1(ram16s_inst_93_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_849 (
  .O(mux_o_849),
  .I0(ram16s_inst_94_dout[1]),
  .I1(ram16s_inst_95_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_850 (
  .O(mux_o_850),
  .I0(ram16s_inst_96_dout[1]),
  .I1(ram16s_inst_97_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_851 (
  .O(mux_o_851),
  .I0(ram16s_inst_98_dout[1]),
  .I1(ram16s_inst_99_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_852 (
  .O(mux_o_852),
  .I0(ram16s_inst_100_dout[1]),
  .I1(ram16s_inst_101_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_853 (
  .O(mux_o_853),
  .I0(ram16s_inst_102_dout[1]),
  .I1(ram16s_inst_103_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_854 (
  .O(mux_o_854),
  .I0(ram16s_inst_104_dout[1]),
  .I1(ram16s_inst_105_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_855 (
  .O(mux_o_855),
  .I0(ram16s_inst_106_dout[1]),
  .I1(ram16s_inst_107_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_856 (
  .O(mux_o_856),
  .I0(ram16s_inst_108_dout[1]),
  .I1(ram16s_inst_109_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_857 (
  .O(mux_o_857),
  .I0(ram16s_inst_110_dout[1]),
  .I1(ram16s_inst_111_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_858 (
  .O(mux_o_858),
  .I0(ram16s_inst_112_dout[1]),
  .I1(ram16s_inst_113_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_859 (
  .O(mux_o_859),
  .I0(ram16s_inst_114_dout[1]),
  .I1(ram16s_inst_115_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_860 (
  .O(mux_o_860),
  .I0(ram16s_inst_116_dout[1]),
  .I1(ram16s_inst_117_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_861 (
  .O(mux_o_861),
  .I0(ram16s_inst_118_dout[1]),
  .I1(ram16s_inst_119_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_862 (
  .O(mux_o_862),
  .I0(ram16s_inst_120_dout[1]),
  .I1(ram16s_inst_121_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_863 (
  .O(mux_o_863),
  .I0(ram16s_inst_122_dout[1]),
  .I1(ram16s_inst_123_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_864 (
  .O(mux_o_864),
  .I0(ram16s_inst_124_dout[1]),
  .I1(ram16s_inst_125_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_865 (
  .O(mux_o_865),
  .I0(ram16s_inst_126_dout[1]),
  .I1(ram16s_inst_127_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_866 (
  .O(mux_o_866),
  .I0(ram16s_inst_128_dout[1]),
  .I1(ram16s_inst_129_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_867 (
  .O(mux_o_867),
  .I0(ram16s_inst_130_dout[1]),
  .I1(ram16s_inst_131_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_868 (
  .O(mux_o_868),
  .I0(ram16s_inst_132_dout[1]),
  .I1(ram16s_inst_133_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_869 (
  .O(mux_o_869),
  .I0(ram16s_inst_134_dout[1]),
  .I1(ram16s_inst_135_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_870 (
  .O(mux_o_870),
  .I0(ram16s_inst_136_dout[1]),
  .I1(ram16s_inst_137_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_871 (
  .O(mux_o_871),
  .I0(ram16s_inst_138_dout[1]),
  .I1(ram16s_inst_139_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_872 (
  .O(mux_o_872),
  .I0(ram16s_inst_140_dout[1]),
  .I1(ram16s_inst_141_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_873 (
  .O(mux_o_873),
  .I0(ram16s_inst_142_dout[1]),
  .I1(ram16s_inst_143_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_874 (
  .O(mux_o_874),
  .I0(ram16s_inst_144_dout[1]),
  .I1(ram16s_inst_145_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_875 (
  .O(mux_o_875),
  .I0(ram16s_inst_146_dout[1]),
  .I1(ram16s_inst_147_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_876 (
  .O(mux_o_876),
  .I0(ram16s_inst_148_dout[1]),
  .I1(ram16s_inst_149_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_877 (
  .O(mux_o_877),
  .I0(ram16s_inst_150_dout[1]),
  .I1(ram16s_inst_151_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_878 (
  .O(mux_o_878),
  .I0(ram16s_inst_152_dout[1]),
  .I1(ram16s_inst_153_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_879 (
  .O(mux_o_879),
  .I0(ram16s_inst_154_dout[1]),
  .I1(ram16s_inst_155_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_880 (
  .O(mux_o_880),
  .I0(ram16s_inst_156_dout[1]),
  .I1(ram16s_inst_157_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_881 (
  .O(mux_o_881),
  .I0(ram16s_inst_158_dout[1]),
  .I1(ram16s_inst_159_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_882 (
  .O(mux_o_882),
  .I0(ram16s_inst_160_dout[1]),
  .I1(ram16s_inst_161_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_883 (
  .O(mux_o_883),
  .I0(ram16s_inst_162_dout[1]),
  .I1(ram16s_inst_163_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_884 (
  .O(mux_o_884),
  .I0(ram16s_inst_164_dout[1]),
  .I1(ram16s_inst_165_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_885 (
  .O(mux_o_885),
  .I0(ram16s_inst_166_dout[1]),
  .I1(ram16s_inst_167_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_886 (
  .O(mux_o_886),
  .I0(ram16s_inst_168_dout[1]),
  .I1(ram16s_inst_169_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_887 (
  .O(mux_o_887),
  .I0(ram16s_inst_170_dout[1]),
  .I1(ram16s_inst_171_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_888 (
  .O(mux_o_888),
  .I0(ram16s_inst_172_dout[1]),
  .I1(ram16s_inst_173_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_889 (
  .O(mux_o_889),
  .I0(ram16s_inst_174_dout[1]),
  .I1(ram16s_inst_175_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_890 (
  .O(mux_o_890),
  .I0(ram16s_inst_176_dout[1]),
  .I1(ram16s_inst_177_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_891 (
  .O(mux_o_891),
  .I0(ram16s_inst_178_dout[1]),
  .I1(ram16s_inst_179_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_892 (
  .O(mux_o_892),
  .I0(ram16s_inst_180_dout[1]),
  .I1(ram16s_inst_181_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_893 (
  .O(mux_o_893),
  .I0(ram16s_inst_182_dout[1]),
  .I1(ram16s_inst_183_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_894 (
  .O(mux_o_894),
  .I0(ram16s_inst_184_dout[1]),
  .I1(ram16s_inst_185_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_895 (
  .O(mux_o_895),
  .I0(ram16s_inst_186_dout[1]),
  .I1(ram16s_inst_187_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_896 (
  .O(mux_o_896),
  .I0(ram16s_inst_188_dout[1]),
  .I1(ram16s_inst_189_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_897 (
  .O(mux_o_897),
  .I0(ram16s_inst_190_dout[1]),
  .I1(ram16s_inst_191_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_898 (
  .O(mux_o_898),
  .I0(ram16s_inst_192_dout[1]),
  .I1(ram16s_inst_193_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_899 (
  .O(mux_o_899),
  .I0(ram16s_inst_194_dout[1]),
  .I1(ram16s_inst_195_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_900 (
  .O(mux_o_900),
  .I0(ram16s_inst_196_dout[1]),
  .I1(ram16s_inst_197_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_901 (
  .O(mux_o_901),
  .I0(ram16s_inst_198_dout[1]),
  .I1(ram16s_inst_199_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_902 (
  .O(mux_o_902),
  .I0(ram16s_inst_200_dout[1]),
  .I1(ram16s_inst_201_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_903 (
  .O(mux_o_903),
  .I0(ram16s_inst_202_dout[1]),
  .I1(ram16s_inst_203_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_904 (
  .O(mux_o_904),
  .I0(ram16s_inst_204_dout[1]),
  .I1(ram16s_inst_205_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_905 (
  .O(mux_o_905),
  .I0(ram16s_inst_206_dout[1]),
  .I1(ram16s_inst_207_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_906 (
  .O(mux_o_906),
  .I0(ram16s_inst_208_dout[1]),
  .I1(ram16s_inst_209_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_907 (
  .O(mux_o_907),
  .I0(ram16s_inst_210_dout[1]),
  .I1(ram16s_inst_211_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_908 (
  .O(mux_o_908),
  .I0(ram16s_inst_212_dout[1]),
  .I1(ram16s_inst_213_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_909 (
  .O(mux_o_909),
  .I0(ram16s_inst_214_dout[1]),
  .I1(ram16s_inst_215_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_910 (
  .O(mux_o_910),
  .I0(ram16s_inst_216_dout[1]),
  .I1(ram16s_inst_217_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_911 (
  .O(mux_o_911),
  .I0(ram16s_inst_218_dout[1]),
  .I1(ram16s_inst_219_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_912 (
  .O(mux_o_912),
  .I0(ram16s_inst_220_dout[1]),
  .I1(ram16s_inst_221_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_913 (
  .O(mux_o_913),
  .I0(ram16s_inst_222_dout[1]),
  .I1(ram16s_inst_223_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_914 (
  .O(mux_o_914),
  .I0(ram16s_inst_224_dout[1]),
  .I1(ram16s_inst_225_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_915 (
  .O(mux_o_915),
  .I0(ram16s_inst_226_dout[1]),
  .I1(ram16s_inst_227_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_916 (
  .O(mux_o_916),
  .I0(ram16s_inst_228_dout[1]),
  .I1(ram16s_inst_229_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_917 (
  .O(mux_o_917),
  .I0(ram16s_inst_230_dout[1]),
  .I1(ram16s_inst_231_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_918 (
  .O(mux_o_918),
  .I0(ram16s_inst_232_dout[1]),
  .I1(ram16s_inst_233_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_919 (
  .O(mux_o_919),
  .I0(ram16s_inst_234_dout[1]),
  .I1(ram16s_inst_235_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_920 (
  .O(mux_o_920),
  .I0(ram16s_inst_236_dout[1]),
  .I1(ram16s_inst_237_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_921 (
  .O(mux_o_921),
  .I0(ram16s_inst_238_dout[1]),
  .I1(ram16s_inst_239_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_922 (
  .O(mux_o_922),
  .I0(ram16s_inst_240_dout[1]),
  .I1(ram16s_inst_241_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_923 (
  .O(mux_o_923),
  .I0(ram16s_inst_242_dout[1]),
  .I1(ram16s_inst_243_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_924 (
  .O(mux_o_924),
  .I0(ram16s_inst_244_dout[1]),
  .I1(ram16s_inst_245_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_925 (
  .O(mux_o_925),
  .I0(ram16s_inst_246_dout[1]),
  .I1(ram16s_inst_247_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_926 (
  .O(mux_o_926),
  .I0(ram16s_inst_248_dout[1]),
  .I1(ram16s_inst_249_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_927 (
  .O(mux_o_927),
  .I0(ram16s_inst_250_dout[1]),
  .I1(ram16s_inst_251_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_928 (
  .O(mux_o_928),
  .I0(ram16s_inst_252_dout[1]),
  .I1(ram16s_inst_253_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_929 (
  .O(mux_o_929),
  .I0(ram16s_inst_254_dout[1]),
  .I1(ram16s_inst_255_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_930 (
  .O(mux_o_930),
  .I0(ram16s_inst_256_dout[1]),
  .I1(ram16s_inst_257_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_931 (
  .O(mux_o_931),
  .I0(ram16s_inst_258_dout[1]),
  .I1(ram16s_inst_259_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_932 (
  .O(mux_o_932),
  .I0(ram16s_inst_260_dout[1]),
  .I1(ram16s_inst_261_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_933 (
  .O(mux_o_933),
  .I0(ram16s_inst_262_dout[1]),
  .I1(ram16s_inst_263_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_934 (
  .O(mux_o_934),
  .I0(ram16s_inst_264_dout[1]),
  .I1(ram16s_inst_265_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_935 (
  .O(mux_o_935),
  .I0(ram16s_inst_266_dout[1]),
  .I1(ram16s_inst_267_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_936 (
  .O(mux_o_936),
  .I0(ram16s_inst_268_dout[1]),
  .I1(ram16s_inst_269_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_937 (
  .O(mux_o_937),
  .I0(ram16s_inst_270_dout[1]),
  .I1(ram16s_inst_271_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_938 (
  .O(mux_o_938),
  .I0(ram16s_inst_272_dout[1]),
  .I1(ram16s_inst_273_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_939 (
  .O(mux_o_939),
  .I0(ram16s_inst_274_dout[1]),
  .I1(ram16s_inst_275_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_940 (
  .O(mux_o_940),
  .I0(ram16s_inst_276_dout[1]),
  .I1(ram16s_inst_277_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_941 (
  .O(mux_o_941),
  .I0(ram16s_inst_278_dout[1]),
  .I1(ram16s_inst_279_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_942 (
  .O(mux_o_942),
  .I0(ram16s_inst_280_dout[1]),
  .I1(ram16s_inst_281_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_943 (
  .O(mux_o_943),
  .I0(ram16s_inst_282_dout[1]),
  .I1(ram16s_inst_283_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_944 (
  .O(mux_o_944),
  .I0(ram16s_inst_284_dout[1]),
  .I1(ram16s_inst_285_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_945 (
  .O(mux_o_945),
  .I0(ram16s_inst_286_dout[1]),
  .I1(ram16s_inst_287_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_946 (
  .O(mux_o_946),
  .I0(ram16s_inst_288_dout[1]),
  .I1(ram16s_inst_289_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_947 (
  .O(mux_o_947),
  .I0(ram16s_inst_290_dout[1]),
  .I1(ram16s_inst_291_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_948 (
  .O(mux_o_948),
  .I0(ram16s_inst_292_dout[1]),
  .I1(ram16s_inst_293_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_949 (
  .O(mux_o_949),
  .I0(ram16s_inst_294_dout[1]),
  .I1(ram16s_inst_295_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_950 (
  .O(mux_o_950),
  .I0(ram16s_inst_296_dout[1]),
  .I1(ram16s_inst_297_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_951 (
  .O(mux_o_951),
  .I0(ram16s_inst_298_dout[1]),
  .I1(ram16s_inst_299_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_952 (
  .O(mux_o_952),
  .I0(ram16s_inst_300_dout[1]),
  .I1(ram16s_inst_301_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_953 (
  .O(mux_o_953),
  .I0(ram16s_inst_302_dout[1]),
  .I1(ram16s_inst_303_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_954 (
  .O(mux_o_954),
  .I0(ram16s_inst_304_dout[1]),
  .I1(ram16s_inst_305_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_955 (
  .O(mux_o_955),
  .I0(ram16s_inst_306_dout[1]),
  .I1(ram16s_inst_307_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_956 (
  .O(mux_o_956),
  .I0(ram16s_inst_308_dout[1]),
  .I1(ram16s_inst_309_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_957 (
  .O(mux_o_957),
  .I0(ram16s_inst_310_dout[1]),
  .I1(ram16s_inst_311_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_958 (
  .O(mux_o_958),
  .I0(ram16s_inst_312_dout[1]),
  .I1(ram16s_inst_313_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_959 (
  .O(mux_o_959),
  .I0(ram16s_inst_314_dout[1]),
  .I1(ram16s_inst_315_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_960 (
  .O(mux_o_960),
  .I0(ram16s_inst_316_dout[1]),
  .I1(ram16s_inst_317_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_961 (
  .O(mux_o_961),
  .I0(ram16s_inst_318_dout[1]),
  .I1(ram16s_inst_319_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_962 (
  .O(mux_o_962),
  .I0(ram16s_inst_320_dout[1]),
  .I1(ram16s_inst_321_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_963 (
  .O(mux_o_963),
  .I0(ram16s_inst_322_dout[1]),
  .I1(ram16s_inst_323_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_964 (
  .O(mux_o_964),
  .I0(ram16s_inst_324_dout[1]),
  .I1(ram16s_inst_325_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_965 (
  .O(mux_o_965),
  .I0(ram16s_inst_326_dout[1]),
  .I1(ram16s_inst_327_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_966 (
  .O(mux_o_966),
  .I0(ram16s_inst_328_dout[1]),
  .I1(ram16s_inst_329_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_967 (
  .O(mux_o_967),
  .I0(ram16s_inst_330_dout[1]),
  .I1(ram16s_inst_331_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_968 (
  .O(mux_o_968),
  .I0(ram16s_inst_332_dout[1]),
  .I1(ram16s_inst_333_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_969 (
  .O(mux_o_969),
  .I0(ram16s_inst_334_dout[1]),
  .I1(ram16s_inst_335_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_970 (
  .O(mux_o_970),
  .I0(ram16s_inst_336_dout[1]),
  .I1(ram16s_inst_337_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_971 (
  .O(mux_o_971),
  .I0(ram16s_inst_338_dout[1]),
  .I1(ram16s_inst_339_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_972 (
  .O(mux_o_972),
  .I0(ram16s_inst_340_dout[1]),
  .I1(ram16s_inst_341_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_973 (
  .O(mux_o_973),
  .I0(ram16s_inst_342_dout[1]),
  .I1(ram16s_inst_343_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_974 (
  .O(mux_o_974),
  .I0(ram16s_inst_344_dout[1]),
  .I1(ram16s_inst_345_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_975 (
  .O(mux_o_975),
  .I0(ram16s_inst_346_dout[1]),
  .I1(ram16s_inst_347_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_976 (
  .O(mux_o_976),
  .I0(ram16s_inst_348_dout[1]),
  .I1(ram16s_inst_349_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_977 (
  .O(mux_o_977),
  .I0(ram16s_inst_350_dout[1]),
  .I1(ram16s_inst_351_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_978 (
  .O(mux_o_978),
  .I0(ram16s_inst_352_dout[1]),
  .I1(ram16s_inst_353_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_979 (
  .O(mux_o_979),
  .I0(ram16s_inst_354_dout[1]),
  .I1(ram16s_inst_355_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_980 (
  .O(mux_o_980),
  .I0(ram16s_inst_356_dout[1]),
  .I1(ram16s_inst_357_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_981 (
  .O(mux_o_981),
  .I0(ram16s_inst_358_dout[1]),
  .I1(ram16s_inst_359_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_982 (
  .O(mux_o_982),
  .I0(ram16s_inst_360_dout[1]),
  .I1(ram16s_inst_361_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_983 (
  .O(mux_o_983),
  .I0(ram16s_inst_362_dout[1]),
  .I1(ram16s_inst_363_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_984 (
  .O(mux_o_984),
  .I0(ram16s_inst_364_dout[1]),
  .I1(ram16s_inst_365_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_985 (
  .O(mux_o_985),
  .I0(ram16s_inst_366_dout[1]),
  .I1(ram16s_inst_367_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_986 (
  .O(mux_o_986),
  .I0(ram16s_inst_368_dout[1]),
  .I1(ram16s_inst_369_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_987 (
  .O(mux_o_987),
  .I0(ram16s_inst_370_dout[1]),
  .I1(ram16s_inst_371_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_988 (
  .O(mux_o_988),
  .I0(ram16s_inst_372_dout[1]),
  .I1(ram16s_inst_373_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_989 (
  .O(mux_o_989),
  .I0(ram16s_inst_374_dout[1]),
  .I1(ram16s_inst_375_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_990 (
  .O(mux_o_990),
  .I0(ram16s_inst_376_dout[1]),
  .I1(ram16s_inst_377_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_991 (
  .O(mux_o_991),
  .I0(ram16s_inst_378_dout[1]),
  .I1(ram16s_inst_379_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_992 (
  .O(mux_o_992),
  .I0(ram16s_inst_380_dout[1]),
  .I1(ram16s_inst_381_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_993 (
  .O(mux_o_993),
  .I0(ram16s_inst_382_dout[1]),
  .I1(ram16s_inst_383_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_994 (
  .O(mux_o_994),
  .I0(ram16s_inst_384_dout[1]),
  .I1(ram16s_inst_385_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_995 (
  .O(mux_o_995),
  .I0(ram16s_inst_386_dout[1]),
  .I1(ram16s_inst_387_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_996 (
  .O(mux_o_996),
  .I0(ram16s_inst_388_dout[1]),
  .I1(ram16s_inst_389_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_997 (
  .O(mux_o_997),
  .I0(ram16s_inst_390_dout[1]),
  .I1(ram16s_inst_391_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_998 (
  .O(mux_o_998),
  .I0(ram16s_inst_392_dout[1]),
  .I1(ram16s_inst_393_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_999 (
  .O(mux_o_999),
  .I0(ram16s_inst_394_dout[1]),
  .I1(ram16s_inst_395_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1000 (
  .O(mux_o_1000),
  .I0(ram16s_inst_396_dout[1]),
  .I1(ram16s_inst_397_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1001 (
  .O(mux_o_1001),
  .I0(ram16s_inst_398_dout[1]),
  .I1(ram16s_inst_399_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1002 (
  .O(mux_o_1002),
  .I0(ram16s_inst_400_dout[1]),
  .I1(ram16s_inst_401_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1003 (
  .O(mux_o_1003),
  .I0(ram16s_inst_402_dout[1]),
  .I1(ram16s_inst_403_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1004 (
  .O(mux_o_1004),
  .I0(ram16s_inst_404_dout[1]),
  .I1(ram16s_inst_405_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1005 (
  .O(mux_o_1005),
  .I0(ram16s_inst_406_dout[1]),
  .I1(ram16s_inst_407_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1006 (
  .O(mux_o_1006),
  .I0(ram16s_inst_408_dout[1]),
  .I1(ram16s_inst_409_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1007 (
  .O(mux_o_1007),
  .I0(ram16s_inst_410_dout[1]),
  .I1(ram16s_inst_411_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1008 (
  .O(mux_o_1008),
  .I0(ram16s_inst_412_dout[1]),
  .I1(ram16s_inst_413_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1009 (
  .O(mux_o_1009),
  .I0(ram16s_inst_414_dout[1]),
  .I1(ram16s_inst_415_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1010 (
  .O(mux_o_1010),
  .I0(ram16s_inst_416_dout[1]),
  .I1(ram16s_inst_417_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1011 (
  .O(mux_o_1011),
  .I0(ram16s_inst_418_dout[1]),
  .I1(ram16s_inst_419_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1012 (
  .O(mux_o_1012),
  .I0(ram16s_inst_420_dout[1]),
  .I1(ram16s_inst_421_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1013 (
  .O(mux_o_1013),
  .I0(ram16s_inst_422_dout[1]),
  .I1(ram16s_inst_423_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1014 (
  .O(mux_o_1014),
  .I0(ram16s_inst_424_dout[1]),
  .I1(ram16s_inst_425_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1015 (
  .O(mux_o_1015),
  .I0(ram16s_inst_426_dout[1]),
  .I1(ram16s_inst_427_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1016 (
  .O(mux_o_1016),
  .I0(ram16s_inst_428_dout[1]),
  .I1(ram16s_inst_429_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1017 (
  .O(mux_o_1017),
  .I0(ram16s_inst_430_dout[1]),
  .I1(ram16s_inst_431_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1018 (
  .O(mux_o_1018),
  .I0(ram16s_inst_432_dout[1]),
  .I1(ram16s_inst_433_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1019 (
  .O(mux_o_1019),
  .I0(ram16s_inst_434_dout[1]),
  .I1(ram16s_inst_435_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1020 (
  .O(mux_o_1020),
  .I0(ram16s_inst_436_dout[1]),
  .I1(ram16s_inst_437_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1021 (
  .O(mux_o_1021),
  .I0(ram16s_inst_438_dout[1]),
  .I1(ram16s_inst_439_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1022 (
  .O(mux_o_1022),
  .I0(ram16s_inst_440_dout[1]),
  .I1(ram16s_inst_441_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1023 (
  .O(mux_o_1023),
  .I0(ram16s_inst_442_dout[1]),
  .I1(ram16s_inst_443_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1024 (
  .O(mux_o_1024),
  .I0(ram16s_inst_444_dout[1]),
  .I1(ram16s_inst_445_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1025 (
  .O(mux_o_1025),
  .I0(ram16s_inst_446_dout[1]),
  .I1(ram16s_inst_447_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1026 (
  .O(mux_o_1026),
  .I0(ram16s_inst_448_dout[1]),
  .I1(ram16s_inst_449_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1027 (
  .O(mux_o_1027),
  .I0(ram16s_inst_450_dout[1]),
  .I1(ram16s_inst_451_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1028 (
  .O(mux_o_1028),
  .I0(ram16s_inst_452_dout[1]),
  .I1(ram16s_inst_453_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1029 (
  .O(mux_o_1029),
  .I0(ram16s_inst_454_dout[1]),
  .I1(ram16s_inst_455_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1030 (
  .O(mux_o_1030),
  .I0(ram16s_inst_456_dout[1]),
  .I1(ram16s_inst_457_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1031 (
  .O(mux_o_1031),
  .I0(ram16s_inst_458_dout[1]),
  .I1(ram16s_inst_459_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1032 (
  .O(mux_o_1032),
  .I0(ram16s_inst_460_dout[1]),
  .I1(ram16s_inst_461_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1033 (
  .O(mux_o_1033),
  .I0(ram16s_inst_462_dout[1]),
  .I1(ram16s_inst_463_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1034 (
  .O(mux_o_1034),
  .I0(ram16s_inst_464_dout[1]),
  .I1(ram16s_inst_465_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1035 (
  .O(mux_o_1035),
  .I0(ram16s_inst_466_dout[1]),
  .I1(ram16s_inst_467_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1036 (
  .O(mux_o_1036),
  .I0(ram16s_inst_468_dout[1]),
  .I1(ram16s_inst_469_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1037 (
  .O(mux_o_1037),
  .I0(ram16s_inst_470_dout[1]),
  .I1(ram16s_inst_471_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1038 (
  .O(mux_o_1038),
  .I0(ram16s_inst_472_dout[1]),
  .I1(ram16s_inst_473_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1039 (
  .O(mux_o_1039),
  .I0(ram16s_inst_474_dout[1]),
  .I1(ram16s_inst_475_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1040 (
  .O(mux_o_1040),
  .I0(ram16s_inst_476_dout[1]),
  .I1(ram16s_inst_477_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1041 (
  .O(mux_o_1041),
  .I0(ram16s_inst_478_dout[1]),
  .I1(ram16s_inst_479_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1042 (
  .O(mux_o_1042),
  .I0(ram16s_inst_480_dout[1]),
  .I1(ram16s_inst_481_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1043 (
  .O(mux_o_1043),
  .I0(ram16s_inst_482_dout[1]),
  .I1(ram16s_inst_483_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1044 (
  .O(mux_o_1044),
  .I0(ram16s_inst_484_dout[1]),
  .I1(ram16s_inst_485_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1045 (
  .O(mux_o_1045),
  .I0(ram16s_inst_486_dout[1]),
  .I1(ram16s_inst_487_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1046 (
  .O(mux_o_1046),
  .I0(ram16s_inst_488_dout[1]),
  .I1(ram16s_inst_489_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1047 (
  .O(mux_o_1047),
  .I0(ram16s_inst_490_dout[1]),
  .I1(ram16s_inst_491_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1048 (
  .O(mux_o_1048),
  .I0(ram16s_inst_492_dout[1]),
  .I1(ram16s_inst_493_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1049 (
  .O(mux_o_1049),
  .I0(ram16s_inst_494_dout[1]),
  .I1(ram16s_inst_495_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1050 (
  .O(mux_o_1050),
  .I0(ram16s_inst_496_dout[1]),
  .I1(ram16s_inst_497_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1051 (
  .O(mux_o_1051),
  .I0(ram16s_inst_498_dout[1]),
  .I1(ram16s_inst_499_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1052 (
  .O(mux_o_1052),
  .I0(ram16s_inst_500_dout[1]),
  .I1(ram16s_inst_501_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1053 (
  .O(mux_o_1053),
  .I0(ram16s_inst_502_dout[1]),
  .I1(ram16s_inst_503_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1054 (
  .O(mux_o_1054),
  .I0(ram16s_inst_504_dout[1]),
  .I1(ram16s_inst_505_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1055 (
  .O(mux_o_1055),
  .I0(ram16s_inst_506_dout[1]),
  .I1(ram16s_inst_507_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1056 (
  .O(mux_o_1056),
  .I0(ram16s_inst_508_dout[1]),
  .I1(ram16s_inst_509_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1057 (
  .O(mux_o_1057),
  .I0(ram16s_inst_510_dout[1]),
  .I1(ram16s_inst_511_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1058 (
  .O(mux_o_1058),
  .I0(ram16s_inst_512_dout[1]),
  .I1(ram16s_inst_513_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1059 (
  .O(mux_o_1059),
  .I0(ram16s_inst_514_dout[1]),
  .I1(ram16s_inst_515_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1060 (
  .O(mux_o_1060),
  .I0(ram16s_inst_516_dout[1]),
  .I1(ram16s_inst_517_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1061 (
  .O(mux_o_1061),
  .I0(ram16s_inst_518_dout[1]),
  .I1(ram16s_inst_519_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1062 (
  .O(mux_o_1062),
  .I0(ram16s_inst_520_dout[1]),
  .I1(ram16s_inst_521_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1063 (
  .O(mux_o_1063),
  .I0(ram16s_inst_522_dout[1]),
  .I1(ram16s_inst_523_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1064 (
  .O(mux_o_1064),
  .I0(ram16s_inst_524_dout[1]),
  .I1(ram16s_inst_525_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1065 (
  .O(mux_o_1065),
  .I0(ram16s_inst_526_dout[1]),
  .I1(ram16s_inst_527_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1066 (
  .O(mux_o_1066),
  .I0(ram16s_inst_528_dout[1]),
  .I1(ram16s_inst_529_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1067 (
  .O(mux_o_1067),
  .I0(ram16s_inst_530_dout[1]),
  .I1(ram16s_inst_531_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1068 (
  .O(mux_o_1068),
  .I0(ram16s_inst_532_dout[1]),
  .I1(ram16s_inst_533_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1069 (
  .O(mux_o_1069),
  .I0(ram16s_inst_534_dout[1]),
  .I1(ram16s_inst_535_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1070 (
  .O(mux_o_1070),
  .I0(ram16s_inst_536_dout[1]),
  .I1(ram16s_inst_537_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1071 (
  .O(mux_o_1071),
  .I0(ram16s_inst_538_dout[1]),
  .I1(ram16s_inst_539_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1072 (
  .O(mux_o_1072),
  .I0(ram16s_inst_540_dout[1]),
  .I1(ram16s_inst_541_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1073 (
  .O(mux_o_1073),
  .I0(ram16s_inst_542_dout[1]),
  .I1(ram16s_inst_543_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1074 (
  .O(mux_o_1074),
  .I0(ram16s_inst_544_dout[1]),
  .I1(ram16s_inst_545_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1075 (
  .O(mux_o_1075),
  .I0(ram16s_inst_546_dout[1]),
  .I1(ram16s_inst_547_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1076 (
  .O(mux_o_1076),
  .I0(ram16s_inst_548_dout[1]),
  .I1(ram16s_inst_549_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1077 (
  .O(mux_o_1077),
  .I0(ram16s_inst_550_dout[1]),
  .I1(ram16s_inst_551_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1078 (
  .O(mux_o_1078),
  .I0(ram16s_inst_552_dout[1]),
  .I1(ram16s_inst_553_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1079 (
  .O(mux_o_1079),
  .I0(ram16s_inst_554_dout[1]),
  .I1(ram16s_inst_555_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1080 (
  .O(mux_o_1080),
  .I0(ram16s_inst_556_dout[1]),
  .I1(ram16s_inst_557_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1081 (
  .O(mux_o_1081),
  .I0(ram16s_inst_558_dout[1]),
  .I1(ram16s_inst_559_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1082 (
  .O(mux_o_1082),
  .I0(ram16s_inst_560_dout[1]),
  .I1(ram16s_inst_561_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1083 (
  .O(mux_o_1083),
  .I0(ram16s_inst_562_dout[1]),
  .I1(ram16s_inst_563_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1084 (
  .O(mux_o_1084),
  .I0(ram16s_inst_564_dout[1]),
  .I1(ram16s_inst_565_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1085 (
  .O(mux_o_1085),
  .I0(ram16s_inst_566_dout[1]),
  .I1(ram16s_inst_567_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1086 (
  .O(mux_o_1086),
  .I0(ram16s_inst_568_dout[1]),
  .I1(ram16s_inst_569_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1087 (
  .O(mux_o_1087),
  .I0(ram16s_inst_570_dout[1]),
  .I1(ram16s_inst_571_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1088 (
  .O(mux_o_1088),
  .I0(ram16s_inst_572_dout[1]),
  .I1(ram16s_inst_573_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1089 (
  .O(mux_o_1089),
  .I0(ram16s_inst_574_dout[1]),
  .I1(ram16s_inst_575_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1090 (
  .O(mux_o_1090),
  .I0(ram16s_inst_576_dout[1]),
  .I1(ram16s_inst_577_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1091 (
  .O(mux_o_1091),
  .I0(ram16s_inst_578_dout[1]),
  .I1(ram16s_inst_579_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1092 (
  .O(mux_o_1092),
  .I0(ram16s_inst_580_dout[1]),
  .I1(ram16s_inst_581_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1093 (
  .O(mux_o_1093),
  .I0(ram16s_inst_582_dout[1]),
  .I1(ram16s_inst_583_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1094 (
  .O(mux_o_1094),
  .I0(ram16s_inst_584_dout[1]),
  .I1(ram16s_inst_585_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1095 (
  .O(mux_o_1095),
  .I0(ram16s_inst_586_dout[1]),
  .I1(ram16s_inst_587_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1096 (
  .O(mux_o_1096),
  .I0(ram16s_inst_588_dout[1]),
  .I1(ram16s_inst_589_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1097 (
  .O(mux_o_1097),
  .I0(ram16s_inst_590_dout[1]),
  .I1(ram16s_inst_591_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1098 (
  .O(mux_o_1098),
  .I0(ram16s_inst_592_dout[1]),
  .I1(ram16s_inst_593_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1099 (
  .O(mux_o_1099),
  .I0(ram16s_inst_594_dout[1]),
  .I1(ram16s_inst_595_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1100 (
  .O(mux_o_1100),
  .I0(ram16s_inst_596_dout[1]),
  .I1(ram16s_inst_597_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1101 (
  .O(mux_o_1101),
  .I0(ram16s_inst_598_dout[1]),
  .I1(ram16s_inst_599_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1102 (
  .O(mux_o_1102),
  .I0(ram16s_inst_600_dout[1]),
  .I1(ram16s_inst_601_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1103 (
  .O(mux_o_1103),
  .I0(ram16s_inst_602_dout[1]),
  .I1(ram16s_inst_603_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1104 (
  .O(mux_o_1104),
  .I0(ram16s_inst_604_dout[1]),
  .I1(ram16s_inst_605_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1105 (
  .O(mux_o_1105),
  .I0(ram16s_inst_606_dout[1]),
  .I1(ram16s_inst_607_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1106 (
  .O(mux_o_1106),
  .I0(ram16s_inst_608_dout[1]),
  .I1(ram16s_inst_609_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1107 (
  .O(mux_o_1107),
  .I0(ram16s_inst_610_dout[1]),
  .I1(ram16s_inst_611_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1108 (
  .O(mux_o_1108),
  .I0(ram16s_inst_612_dout[1]),
  .I1(ram16s_inst_613_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1109 (
  .O(mux_o_1109),
  .I0(ram16s_inst_614_dout[1]),
  .I1(ram16s_inst_615_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1110 (
  .O(mux_o_1110),
  .I0(ram16s_inst_616_dout[1]),
  .I1(ram16s_inst_617_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1111 (
  .O(mux_o_1111),
  .I0(ram16s_inst_618_dout[1]),
  .I1(ram16s_inst_619_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1112 (
  .O(mux_o_1112),
  .I0(ram16s_inst_620_dout[1]),
  .I1(ram16s_inst_621_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1113 (
  .O(mux_o_1113),
  .I0(ram16s_inst_622_dout[1]),
  .I1(ram16s_inst_623_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1114 (
  .O(mux_o_1114),
  .I0(ram16s_inst_624_dout[1]),
  .I1(ram16s_inst_625_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1115 (
  .O(mux_o_1115),
  .I0(ram16s_inst_626_dout[1]),
  .I1(ram16s_inst_627_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1116 (
  .O(mux_o_1116),
  .I0(ram16s_inst_628_dout[1]),
  .I1(ram16s_inst_629_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1117 (
  .O(mux_o_1117),
  .I0(ram16s_inst_630_dout[1]),
  .I1(ram16s_inst_631_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1118 (
  .O(mux_o_1118),
  .I0(ram16s_inst_632_dout[1]),
  .I1(ram16s_inst_633_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1119 (
  .O(mux_o_1119),
  .I0(ram16s_inst_634_dout[1]),
  .I1(ram16s_inst_635_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1120 (
  .O(mux_o_1120),
  .I0(ram16s_inst_636_dout[1]),
  .I1(ram16s_inst_637_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1121 (
  .O(mux_o_1121),
  .I0(ram16s_inst_638_dout[1]),
  .I1(ram16s_inst_639_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1122 (
  .O(mux_o_1122),
  .I0(ram16s_inst_640_dout[1]),
  .I1(ram16s_inst_641_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1123 (
  .O(mux_o_1123),
  .I0(ram16s_inst_642_dout[1]),
  .I1(ram16s_inst_643_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1124 (
  .O(mux_o_1124),
  .I0(ram16s_inst_644_dout[1]),
  .I1(ram16s_inst_645_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1125 (
  .O(mux_o_1125),
  .I0(ram16s_inst_646_dout[1]),
  .I1(ram16s_inst_647_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1126 (
  .O(mux_o_1126),
  .I0(ram16s_inst_648_dout[1]),
  .I1(ram16s_inst_649_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1127 (
  .O(mux_o_1127),
  .I0(ram16s_inst_650_dout[1]),
  .I1(ram16s_inst_651_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1128 (
  .O(mux_o_1128),
  .I0(ram16s_inst_652_dout[1]),
  .I1(ram16s_inst_653_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1129 (
  .O(mux_o_1129),
  .I0(ram16s_inst_654_dout[1]),
  .I1(ram16s_inst_655_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1130 (
  .O(mux_o_1130),
  .I0(ram16s_inst_656_dout[1]),
  .I1(ram16s_inst_657_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1131 (
  .O(mux_o_1131),
  .I0(ram16s_inst_658_dout[1]),
  .I1(ram16s_inst_659_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1132 (
  .O(mux_o_1132),
  .I0(ram16s_inst_660_dout[1]),
  .I1(ram16s_inst_661_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1133 (
  .O(mux_o_1133),
  .I0(ram16s_inst_662_dout[1]),
  .I1(ram16s_inst_663_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1134 (
  .O(mux_o_1134),
  .I0(ram16s_inst_664_dout[1]),
  .I1(ram16s_inst_665_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1135 (
  .O(mux_o_1135),
  .I0(ram16s_inst_666_dout[1]),
  .I1(ram16s_inst_667_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1136 (
  .O(mux_o_1136),
  .I0(ram16s_inst_668_dout[1]),
  .I1(ram16s_inst_669_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1137 (
  .O(mux_o_1137),
  .I0(ram16s_inst_670_dout[1]),
  .I1(ram16s_inst_671_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1138 (
  .O(mux_o_1138),
  .I0(ram16s_inst_672_dout[1]),
  .I1(ram16s_inst_673_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1139 (
  .O(mux_o_1139),
  .I0(ram16s_inst_674_dout[1]),
  .I1(ram16s_inst_675_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1140 (
  .O(mux_o_1140),
  .I0(ram16s_inst_676_dout[1]),
  .I1(ram16s_inst_677_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1141 (
  .O(mux_o_1141),
  .I0(ram16s_inst_678_dout[1]),
  .I1(ram16s_inst_679_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1142 (
  .O(mux_o_1142),
  .I0(ram16s_inst_680_dout[1]),
  .I1(ram16s_inst_681_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1143 (
  .O(mux_o_1143),
  .I0(ram16s_inst_682_dout[1]),
  .I1(ram16s_inst_683_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1144 (
  .O(mux_o_1144),
  .I0(ram16s_inst_684_dout[1]),
  .I1(ram16s_inst_685_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1145 (
  .O(mux_o_1145),
  .I0(ram16s_inst_686_dout[1]),
  .I1(ram16s_inst_687_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1146 (
  .O(mux_o_1146),
  .I0(ram16s_inst_688_dout[1]),
  .I1(ram16s_inst_689_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1147 (
  .O(mux_o_1147),
  .I0(ram16s_inst_690_dout[1]),
  .I1(ram16s_inst_691_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1148 (
  .O(mux_o_1148),
  .I0(ram16s_inst_692_dout[1]),
  .I1(ram16s_inst_693_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1149 (
  .O(mux_o_1149),
  .I0(ram16s_inst_694_dout[1]),
  .I1(ram16s_inst_695_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1150 (
  .O(mux_o_1150),
  .I0(ram16s_inst_696_dout[1]),
  .I1(ram16s_inst_697_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1151 (
  .O(mux_o_1151),
  .I0(ram16s_inst_698_dout[1]),
  .I1(ram16s_inst_699_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1152 (
  .O(mux_o_1152),
  .I0(ram16s_inst_700_dout[1]),
  .I1(ram16s_inst_701_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1153 (
  .O(mux_o_1153),
  .I0(ram16s_inst_702_dout[1]),
  .I1(ram16s_inst_703_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1154 (
  .O(mux_o_1154),
  .I0(ram16s_inst_704_dout[1]),
  .I1(ram16s_inst_705_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1155 (
  .O(mux_o_1155),
  .I0(ram16s_inst_706_dout[1]),
  .I1(ram16s_inst_707_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1156 (
  .O(mux_o_1156),
  .I0(ram16s_inst_708_dout[1]),
  .I1(ram16s_inst_709_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1157 (
  .O(mux_o_1157),
  .I0(ram16s_inst_710_dout[1]),
  .I1(ram16s_inst_711_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1158 (
  .O(mux_o_1158),
  .I0(ram16s_inst_712_dout[1]),
  .I1(ram16s_inst_713_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1159 (
  .O(mux_o_1159),
  .I0(ram16s_inst_714_dout[1]),
  .I1(ram16s_inst_715_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1160 (
  .O(mux_o_1160),
  .I0(ram16s_inst_716_dout[1]),
  .I1(ram16s_inst_717_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1161 (
  .O(mux_o_1161),
  .I0(ram16s_inst_718_dout[1]),
  .I1(ram16s_inst_719_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1162 (
  .O(mux_o_1162),
  .I0(ram16s_inst_720_dout[1]),
  .I1(ram16s_inst_721_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1163 (
  .O(mux_o_1163),
  .I0(ram16s_inst_722_dout[1]),
  .I1(ram16s_inst_723_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1164 (
  .O(mux_o_1164),
  .I0(ram16s_inst_724_dout[1]),
  .I1(ram16s_inst_725_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1165 (
  .O(mux_o_1165),
  .I0(ram16s_inst_726_dout[1]),
  .I1(ram16s_inst_727_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1166 (
  .O(mux_o_1166),
  .I0(ram16s_inst_728_dout[1]),
  .I1(ram16s_inst_729_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1167 (
  .O(mux_o_1167),
  .I0(ram16s_inst_730_dout[1]),
  .I1(ram16s_inst_731_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1168 (
  .O(mux_o_1168),
  .I0(ram16s_inst_732_dout[1]),
  .I1(ram16s_inst_733_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1169 (
  .O(mux_o_1169),
  .I0(ram16s_inst_734_dout[1]),
  .I1(ram16s_inst_735_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1170 (
  .O(mux_o_1170),
  .I0(ram16s_inst_736_dout[1]),
  .I1(ram16s_inst_737_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1171 (
  .O(mux_o_1171),
  .I0(ram16s_inst_738_dout[1]),
  .I1(ram16s_inst_739_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1172 (
  .O(mux_o_1172),
  .I0(ram16s_inst_740_dout[1]),
  .I1(ram16s_inst_741_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1173 (
  .O(mux_o_1173),
  .I0(ram16s_inst_742_dout[1]),
  .I1(ram16s_inst_743_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1174 (
  .O(mux_o_1174),
  .I0(ram16s_inst_744_dout[1]),
  .I1(ram16s_inst_745_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1175 (
  .O(mux_o_1175),
  .I0(ram16s_inst_746_dout[1]),
  .I1(ram16s_inst_747_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1176 (
  .O(mux_o_1176),
  .I0(ram16s_inst_748_dout[1]),
  .I1(ram16s_inst_749_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1177 (
  .O(mux_o_1177),
  .I0(ram16s_inst_750_dout[1]),
  .I1(ram16s_inst_751_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1178 (
  .O(mux_o_1178),
  .I0(ram16s_inst_752_dout[1]),
  .I1(ram16s_inst_753_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1179 (
  .O(mux_o_1179),
  .I0(ram16s_inst_754_dout[1]),
  .I1(ram16s_inst_755_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1180 (
  .O(mux_o_1180),
  .I0(ram16s_inst_756_dout[1]),
  .I1(ram16s_inst_757_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1181 (
  .O(mux_o_1181),
  .I0(ram16s_inst_758_dout[1]),
  .I1(ram16s_inst_759_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1182 (
  .O(mux_o_1182),
  .I0(ram16s_inst_760_dout[1]),
  .I1(ram16s_inst_761_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1183 (
  .O(mux_o_1183),
  .I0(ram16s_inst_762_dout[1]),
  .I1(ram16s_inst_763_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1184 (
  .O(mux_o_1184),
  .I0(ram16s_inst_764_dout[1]),
  .I1(ram16s_inst_765_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1185 (
  .O(mux_o_1185),
  .I0(ram16s_inst_766_dout[1]),
  .I1(ram16s_inst_767_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1186 (
  .O(mux_o_1186),
  .I0(ram16s_inst_768_dout[1]),
  .I1(ram16s_inst_769_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1187 (
  .O(mux_o_1187),
  .I0(ram16s_inst_770_dout[1]),
  .I1(ram16s_inst_771_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1188 (
  .O(mux_o_1188),
  .I0(ram16s_inst_772_dout[1]),
  .I1(ram16s_inst_773_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1189 (
  .O(mux_o_1189),
  .I0(ram16s_inst_774_dout[1]),
  .I1(ram16s_inst_775_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1190 (
  .O(mux_o_1190),
  .I0(ram16s_inst_776_dout[1]),
  .I1(ram16s_inst_777_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1191 (
  .O(mux_o_1191),
  .I0(ram16s_inst_778_dout[1]),
  .I1(ram16s_inst_779_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1192 (
  .O(mux_o_1192),
  .I0(ram16s_inst_780_dout[1]),
  .I1(ram16s_inst_781_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1193 (
  .O(mux_o_1193),
  .I0(ram16s_inst_782_dout[1]),
  .I1(ram16s_inst_783_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1194 (
  .O(mux_o_1194),
  .I0(ram16s_inst_784_dout[1]),
  .I1(ram16s_inst_785_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1195 (
  .O(mux_o_1195),
  .I0(ram16s_inst_786_dout[1]),
  .I1(ram16s_inst_787_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1196 (
  .O(mux_o_1196),
  .I0(ram16s_inst_788_dout[1]),
  .I1(ram16s_inst_789_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1197 (
  .O(mux_o_1197),
  .I0(ram16s_inst_790_dout[1]),
  .I1(ram16s_inst_791_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1198 (
  .O(mux_o_1198),
  .I0(ram16s_inst_792_dout[1]),
  .I1(ram16s_inst_793_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1199 (
  .O(mux_o_1199),
  .I0(ram16s_inst_794_dout[1]),
  .I1(ram16s_inst_795_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1200 (
  .O(mux_o_1200),
  .I0(ram16s_inst_796_dout[1]),
  .I1(ram16s_inst_797_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1201 (
  .O(mux_o_1201),
  .I0(ram16s_inst_798_dout[1]),
  .I1(ram16s_inst_799_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_1202 (
  .O(mux_o_1202),
  .I0(mux_o_802),
  .I1(mux_o_803),
  .S0(ad[5])
);
MUX2 mux_inst_1203 (
  .O(mux_o_1203),
  .I0(mux_o_804),
  .I1(mux_o_805),
  .S0(ad[5])
);
MUX2 mux_inst_1204 (
  .O(mux_o_1204),
  .I0(mux_o_806),
  .I1(mux_o_807),
  .S0(ad[5])
);
MUX2 mux_inst_1205 (
  .O(mux_o_1205),
  .I0(mux_o_808),
  .I1(mux_o_809),
  .S0(ad[5])
);
MUX2 mux_inst_1206 (
  .O(mux_o_1206),
  .I0(mux_o_810),
  .I1(mux_o_811),
  .S0(ad[5])
);
MUX2 mux_inst_1207 (
  .O(mux_o_1207),
  .I0(mux_o_812),
  .I1(mux_o_813),
  .S0(ad[5])
);
MUX2 mux_inst_1208 (
  .O(mux_o_1208),
  .I0(mux_o_814),
  .I1(mux_o_815),
  .S0(ad[5])
);
MUX2 mux_inst_1209 (
  .O(mux_o_1209),
  .I0(mux_o_816),
  .I1(mux_o_817),
  .S0(ad[5])
);
MUX2 mux_inst_1210 (
  .O(mux_o_1210),
  .I0(mux_o_818),
  .I1(mux_o_819),
  .S0(ad[5])
);
MUX2 mux_inst_1211 (
  .O(mux_o_1211),
  .I0(mux_o_820),
  .I1(mux_o_821),
  .S0(ad[5])
);
MUX2 mux_inst_1212 (
  .O(mux_o_1212),
  .I0(mux_o_822),
  .I1(mux_o_823),
  .S0(ad[5])
);
MUX2 mux_inst_1213 (
  .O(mux_o_1213),
  .I0(mux_o_824),
  .I1(mux_o_825),
  .S0(ad[5])
);
MUX2 mux_inst_1214 (
  .O(mux_o_1214),
  .I0(mux_o_826),
  .I1(mux_o_827),
  .S0(ad[5])
);
MUX2 mux_inst_1215 (
  .O(mux_o_1215),
  .I0(mux_o_828),
  .I1(mux_o_829),
  .S0(ad[5])
);
MUX2 mux_inst_1216 (
  .O(mux_o_1216),
  .I0(mux_o_830),
  .I1(mux_o_831),
  .S0(ad[5])
);
MUX2 mux_inst_1217 (
  .O(mux_o_1217),
  .I0(mux_o_832),
  .I1(mux_o_833),
  .S0(ad[5])
);
MUX2 mux_inst_1218 (
  .O(mux_o_1218),
  .I0(mux_o_834),
  .I1(mux_o_835),
  .S0(ad[5])
);
MUX2 mux_inst_1219 (
  .O(mux_o_1219),
  .I0(mux_o_836),
  .I1(mux_o_837),
  .S0(ad[5])
);
MUX2 mux_inst_1220 (
  .O(mux_o_1220),
  .I0(mux_o_838),
  .I1(mux_o_839),
  .S0(ad[5])
);
MUX2 mux_inst_1221 (
  .O(mux_o_1221),
  .I0(mux_o_840),
  .I1(mux_o_841),
  .S0(ad[5])
);
MUX2 mux_inst_1222 (
  .O(mux_o_1222),
  .I0(mux_o_842),
  .I1(mux_o_843),
  .S0(ad[5])
);
MUX2 mux_inst_1223 (
  .O(mux_o_1223),
  .I0(mux_o_844),
  .I1(mux_o_845),
  .S0(ad[5])
);
MUX2 mux_inst_1224 (
  .O(mux_o_1224),
  .I0(mux_o_846),
  .I1(mux_o_847),
  .S0(ad[5])
);
MUX2 mux_inst_1225 (
  .O(mux_o_1225),
  .I0(mux_o_848),
  .I1(mux_o_849),
  .S0(ad[5])
);
MUX2 mux_inst_1226 (
  .O(mux_o_1226),
  .I0(mux_o_850),
  .I1(mux_o_851),
  .S0(ad[5])
);
MUX2 mux_inst_1227 (
  .O(mux_o_1227),
  .I0(mux_o_852),
  .I1(mux_o_853),
  .S0(ad[5])
);
MUX2 mux_inst_1228 (
  .O(mux_o_1228),
  .I0(mux_o_854),
  .I1(mux_o_855),
  .S0(ad[5])
);
MUX2 mux_inst_1229 (
  .O(mux_o_1229),
  .I0(mux_o_856),
  .I1(mux_o_857),
  .S0(ad[5])
);
MUX2 mux_inst_1230 (
  .O(mux_o_1230),
  .I0(mux_o_858),
  .I1(mux_o_859),
  .S0(ad[5])
);
MUX2 mux_inst_1231 (
  .O(mux_o_1231),
  .I0(mux_o_860),
  .I1(mux_o_861),
  .S0(ad[5])
);
MUX2 mux_inst_1232 (
  .O(mux_o_1232),
  .I0(mux_o_862),
  .I1(mux_o_863),
  .S0(ad[5])
);
MUX2 mux_inst_1233 (
  .O(mux_o_1233),
  .I0(mux_o_864),
  .I1(mux_o_865),
  .S0(ad[5])
);
MUX2 mux_inst_1234 (
  .O(mux_o_1234),
  .I0(mux_o_866),
  .I1(mux_o_867),
  .S0(ad[5])
);
MUX2 mux_inst_1235 (
  .O(mux_o_1235),
  .I0(mux_o_868),
  .I1(mux_o_869),
  .S0(ad[5])
);
MUX2 mux_inst_1236 (
  .O(mux_o_1236),
  .I0(mux_o_870),
  .I1(mux_o_871),
  .S0(ad[5])
);
MUX2 mux_inst_1237 (
  .O(mux_o_1237),
  .I0(mux_o_872),
  .I1(mux_o_873),
  .S0(ad[5])
);
MUX2 mux_inst_1238 (
  .O(mux_o_1238),
  .I0(mux_o_874),
  .I1(mux_o_875),
  .S0(ad[5])
);
MUX2 mux_inst_1239 (
  .O(mux_o_1239),
  .I0(mux_o_876),
  .I1(mux_o_877),
  .S0(ad[5])
);
MUX2 mux_inst_1240 (
  .O(mux_o_1240),
  .I0(mux_o_878),
  .I1(mux_o_879),
  .S0(ad[5])
);
MUX2 mux_inst_1241 (
  .O(mux_o_1241),
  .I0(mux_o_880),
  .I1(mux_o_881),
  .S0(ad[5])
);
MUX2 mux_inst_1242 (
  .O(mux_o_1242),
  .I0(mux_o_882),
  .I1(mux_o_883),
  .S0(ad[5])
);
MUX2 mux_inst_1243 (
  .O(mux_o_1243),
  .I0(mux_o_884),
  .I1(mux_o_885),
  .S0(ad[5])
);
MUX2 mux_inst_1244 (
  .O(mux_o_1244),
  .I0(mux_o_886),
  .I1(mux_o_887),
  .S0(ad[5])
);
MUX2 mux_inst_1245 (
  .O(mux_o_1245),
  .I0(mux_o_888),
  .I1(mux_o_889),
  .S0(ad[5])
);
MUX2 mux_inst_1246 (
  .O(mux_o_1246),
  .I0(mux_o_890),
  .I1(mux_o_891),
  .S0(ad[5])
);
MUX2 mux_inst_1247 (
  .O(mux_o_1247),
  .I0(mux_o_892),
  .I1(mux_o_893),
  .S0(ad[5])
);
MUX2 mux_inst_1248 (
  .O(mux_o_1248),
  .I0(mux_o_894),
  .I1(mux_o_895),
  .S0(ad[5])
);
MUX2 mux_inst_1249 (
  .O(mux_o_1249),
  .I0(mux_o_896),
  .I1(mux_o_897),
  .S0(ad[5])
);
MUX2 mux_inst_1250 (
  .O(mux_o_1250),
  .I0(mux_o_898),
  .I1(mux_o_899),
  .S0(ad[5])
);
MUX2 mux_inst_1251 (
  .O(mux_o_1251),
  .I0(mux_o_900),
  .I1(mux_o_901),
  .S0(ad[5])
);
MUX2 mux_inst_1252 (
  .O(mux_o_1252),
  .I0(mux_o_902),
  .I1(mux_o_903),
  .S0(ad[5])
);
MUX2 mux_inst_1253 (
  .O(mux_o_1253),
  .I0(mux_o_904),
  .I1(mux_o_905),
  .S0(ad[5])
);
MUX2 mux_inst_1254 (
  .O(mux_o_1254),
  .I0(mux_o_906),
  .I1(mux_o_907),
  .S0(ad[5])
);
MUX2 mux_inst_1255 (
  .O(mux_o_1255),
  .I0(mux_o_908),
  .I1(mux_o_909),
  .S0(ad[5])
);
MUX2 mux_inst_1256 (
  .O(mux_o_1256),
  .I0(mux_o_910),
  .I1(mux_o_911),
  .S0(ad[5])
);
MUX2 mux_inst_1257 (
  .O(mux_o_1257),
  .I0(mux_o_912),
  .I1(mux_o_913),
  .S0(ad[5])
);
MUX2 mux_inst_1258 (
  .O(mux_o_1258),
  .I0(mux_o_914),
  .I1(mux_o_915),
  .S0(ad[5])
);
MUX2 mux_inst_1259 (
  .O(mux_o_1259),
  .I0(mux_o_916),
  .I1(mux_o_917),
  .S0(ad[5])
);
MUX2 mux_inst_1260 (
  .O(mux_o_1260),
  .I0(mux_o_918),
  .I1(mux_o_919),
  .S0(ad[5])
);
MUX2 mux_inst_1261 (
  .O(mux_o_1261),
  .I0(mux_o_920),
  .I1(mux_o_921),
  .S0(ad[5])
);
MUX2 mux_inst_1262 (
  .O(mux_o_1262),
  .I0(mux_o_922),
  .I1(mux_o_923),
  .S0(ad[5])
);
MUX2 mux_inst_1263 (
  .O(mux_o_1263),
  .I0(mux_o_924),
  .I1(mux_o_925),
  .S0(ad[5])
);
MUX2 mux_inst_1264 (
  .O(mux_o_1264),
  .I0(mux_o_926),
  .I1(mux_o_927),
  .S0(ad[5])
);
MUX2 mux_inst_1265 (
  .O(mux_o_1265),
  .I0(mux_o_928),
  .I1(mux_o_929),
  .S0(ad[5])
);
MUX2 mux_inst_1266 (
  .O(mux_o_1266),
  .I0(mux_o_930),
  .I1(mux_o_931),
  .S0(ad[5])
);
MUX2 mux_inst_1267 (
  .O(mux_o_1267),
  .I0(mux_o_932),
  .I1(mux_o_933),
  .S0(ad[5])
);
MUX2 mux_inst_1268 (
  .O(mux_o_1268),
  .I0(mux_o_934),
  .I1(mux_o_935),
  .S0(ad[5])
);
MUX2 mux_inst_1269 (
  .O(mux_o_1269),
  .I0(mux_o_936),
  .I1(mux_o_937),
  .S0(ad[5])
);
MUX2 mux_inst_1270 (
  .O(mux_o_1270),
  .I0(mux_o_938),
  .I1(mux_o_939),
  .S0(ad[5])
);
MUX2 mux_inst_1271 (
  .O(mux_o_1271),
  .I0(mux_o_940),
  .I1(mux_o_941),
  .S0(ad[5])
);
MUX2 mux_inst_1272 (
  .O(mux_o_1272),
  .I0(mux_o_942),
  .I1(mux_o_943),
  .S0(ad[5])
);
MUX2 mux_inst_1273 (
  .O(mux_o_1273),
  .I0(mux_o_944),
  .I1(mux_o_945),
  .S0(ad[5])
);
MUX2 mux_inst_1274 (
  .O(mux_o_1274),
  .I0(mux_o_946),
  .I1(mux_o_947),
  .S0(ad[5])
);
MUX2 mux_inst_1275 (
  .O(mux_o_1275),
  .I0(mux_o_948),
  .I1(mux_o_949),
  .S0(ad[5])
);
MUX2 mux_inst_1276 (
  .O(mux_o_1276),
  .I0(mux_o_950),
  .I1(mux_o_951),
  .S0(ad[5])
);
MUX2 mux_inst_1277 (
  .O(mux_o_1277),
  .I0(mux_o_952),
  .I1(mux_o_953),
  .S0(ad[5])
);
MUX2 mux_inst_1278 (
  .O(mux_o_1278),
  .I0(mux_o_954),
  .I1(mux_o_955),
  .S0(ad[5])
);
MUX2 mux_inst_1279 (
  .O(mux_o_1279),
  .I0(mux_o_956),
  .I1(mux_o_957),
  .S0(ad[5])
);
MUX2 mux_inst_1280 (
  .O(mux_o_1280),
  .I0(mux_o_958),
  .I1(mux_o_959),
  .S0(ad[5])
);
MUX2 mux_inst_1281 (
  .O(mux_o_1281),
  .I0(mux_o_960),
  .I1(mux_o_961),
  .S0(ad[5])
);
MUX2 mux_inst_1282 (
  .O(mux_o_1282),
  .I0(mux_o_962),
  .I1(mux_o_963),
  .S0(ad[5])
);
MUX2 mux_inst_1283 (
  .O(mux_o_1283),
  .I0(mux_o_964),
  .I1(mux_o_965),
  .S0(ad[5])
);
MUX2 mux_inst_1284 (
  .O(mux_o_1284),
  .I0(mux_o_966),
  .I1(mux_o_967),
  .S0(ad[5])
);
MUX2 mux_inst_1285 (
  .O(mux_o_1285),
  .I0(mux_o_968),
  .I1(mux_o_969),
  .S0(ad[5])
);
MUX2 mux_inst_1286 (
  .O(mux_o_1286),
  .I0(mux_o_970),
  .I1(mux_o_971),
  .S0(ad[5])
);
MUX2 mux_inst_1287 (
  .O(mux_o_1287),
  .I0(mux_o_972),
  .I1(mux_o_973),
  .S0(ad[5])
);
MUX2 mux_inst_1288 (
  .O(mux_o_1288),
  .I0(mux_o_974),
  .I1(mux_o_975),
  .S0(ad[5])
);
MUX2 mux_inst_1289 (
  .O(mux_o_1289),
  .I0(mux_o_976),
  .I1(mux_o_977),
  .S0(ad[5])
);
MUX2 mux_inst_1290 (
  .O(mux_o_1290),
  .I0(mux_o_978),
  .I1(mux_o_979),
  .S0(ad[5])
);
MUX2 mux_inst_1291 (
  .O(mux_o_1291),
  .I0(mux_o_980),
  .I1(mux_o_981),
  .S0(ad[5])
);
MUX2 mux_inst_1292 (
  .O(mux_o_1292),
  .I0(mux_o_982),
  .I1(mux_o_983),
  .S0(ad[5])
);
MUX2 mux_inst_1293 (
  .O(mux_o_1293),
  .I0(mux_o_984),
  .I1(mux_o_985),
  .S0(ad[5])
);
MUX2 mux_inst_1294 (
  .O(mux_o_1294),
  .I0(mux_o_986),
  .I1(mux_o_987),
  .S0(ad[5])
);
MUX2 mux_inst_1295 (
  .O(mux_o_1295),
  .I0(mux_o_988),
  .I1(mux_o_989),
  .S0(ad[5])
);
MUX2 mux_inst_1296 (
  .O(mux_o_1296),
  .I0(mux_o_990),
  .I1(mux_o_991),
  .S0(ad[5])
);
MUX2 mux_inst_1297 (
  .O(mux_o_1297),
  .I0(mux_o_992),
  .I1(mux_o_993),
  .S0(ad[5])
);
MUX2 mux_inst_1298 (
  .O(mux_o_1298),
  .I0(mux_o_994),
  .I1(mux_o_995),
  .S0(ad[5])
);
MUX2 mux_inst_1299 (
  .O(mux_o_1299),
  .I0(mux_o_996),
  .I1(mux_o_997),
  .S0(ad[5])
);
MUX2 mux_inst_1300 (
  .O(mux_o_1300),
  .I0(mux_o_998),
  .I1(mux_o_999),
  .S0(ad[5])
);
MUX2 mux_inst_1301 (
  .O(mux_o_1301),
  .I0(mux_o_1000),
  .I1(mux_o_1001),
  .S0(ad[5])
);
MUX2 mux_inst_1302 (
  .O(mux_o_1302),
  .I0(mux_o_1002),
  .I1(mux_o_1003),
  .S0(ad[5])
);
MUX2 mux_inst_1303 (
  .O(mux_o_1303),
  .I0(mux_o_1004),
  .I1(mux_o_1005),
  .S0(ad[5])
);
MUX2 mux_inst_1304 (
  .O(mux_o_1304),
  .I0(mux_o_1006),
  .I1(mux_o_1007),
  .S0(ad[5])
);
MUX2 mux_inst_1305 (
  .O(mux_o_1305),
  .I0(mux_o_1008),
  .I1(mux_o_1009),
  .S0(ad[5])
);
MUX2 mux_inst_1306 (
  .O(mux_o_1306),
  .I0(mux_o_1010),
  .I1(mux_o_1011),
  .S0(ad[5])
);
MUX2 mux_inst_1307 (
  .O(mux_o_1307),
  .I0(mux_o_1012),
  .I1(mux_o_1013),
  .S0(ad[5])
);
MUX2 mux_inst_1308 (
  .O(mux_o_1308),
  .I0(mux_o_1014),
  .I1(mux_o_1015),
  .S0(ad[5])
);
MUX2 mux_inst_1309 (
  .O(mux_o_1309),
  .I0(mux_o_1016),
  .I1(mux_o_1017),
  .S0(ad[5])
);
MUX2 mux_inst_1310 (
  .O(mux_o_1310),
  .I0(mux_o_1018),
  .I1(mux_o_1019),
  .S0(ad[5])
);
MUX2 mux_inst_1311 (
  .O(mux_o_1311),
  .I0(mux_o_1020),
  .I1(mux_o_1021),
  .S0(ad[5])
);
MUX2 mux_inst_1312 (
  .O(mux_o_1312),
  .I0(mux_o_1022),
  .I1(mux_o_1023),
  .S0(ad[5])
);
MUX2 mux_inst_1313 (
  .O(mux_o_1313),
  .I0(mux_o_1024),
  .I1(mux_o_1025),
  .S0(ad[5])
);
MUX2 mux_inst_1314 (
  .O(mux_o_1314),
  .I0(mux_o_1026),
  .I1(mux_o_1027),
  .S0(ad[5])
);
MUX2 mux_inst_1315 (
  .O(mux_o_1315),
  .I0(mux_o_1028),
  .I1(mux_o_1029),
  .S0(ad[5])
);
MUX2 mux_inst_1316 (
  .O(mux_o_1316),
  .I0(mux_o_1030),
  .I1(mux_o_1031),
  .S0(ad[5])
);
MUX2 mux_inst_1317 (
  .O(mux_o_1317),
  .I0(mux_o_1032),
  .I1(mux_o_1033),
  .S0(ad[5])
);
MUX2 mux_inst_1318 (
  .O(mux_o_1318),
  .I0(mux_o_1034),
  .I1(mux_o_1035),
  .S0(ad[5])
);
MUX2 mux_inst_1319 (
  .O(mux_o_1319),
  .I0(mux_o_1036),
  .I1(mux_o_1037),
  .S0(ad[5])
);
MUX2 mux_inst_1320 (
  .O(mux_o_1320),
  .I0(mux_o_1038),
  .I1(mux_o_1039),
  .S0(ad[5])
);
MUX2 mux_inst_1321 (
  .O(mux_o_1321),
  .I0(mux_o_1040),
  .I1(mux_o_1041),
  .S0(ad[5])
);
MUX2 mux_inst_1322 (
  .O(mux_o_1322),
  .I0(mux_o_1042),
  .I1(mux_o_1043),
  .S0(ad[5])
);
MUX2 mux_inst_1323 (
  .O(mux_o_1323),
  .I0(mux_o_1044),
  .I1(mux_o_1045),
  .S0(ad[5])
);
MUX2 mux_inst_1324 (
  .O(mux_o_1324),
  .I0(mux_o_1046),
  .I1(mux_o_1047),
  .S0(ad[5])
);
MUX2 mux_inst_1325 (
  .O(mux_o_1325),
  .I0(mux_o_1048),
  .I1(mux_o_1049),
  .S0(ad[5])
);
MUX2 mux_inst_1326 (
  .O(mux_o_1326),
  .I0(mux_o_1050),
  .I1(mux_o_1051),
  .S0(ad[5])
);
MUX2 mux_inst_1327 (
  .O(mux_o_1327),
  .I0(mux_o_1052),
  .I1(mux_o_1053),
  .S0(ad[5])
);
MUX2 mux_inst_1328 (
  .O(mux_o_1328),
  .I0(mux_o_1054),
  .I1(mux_o_1055),
  .S0(ad[5])
);
MUX2 mux_inst_1329 (
  .O(mux_o_1329),
  .I0(mux_o_1056),
  .I1(mux_o_1057),
  .S0(ad[5])
);
MUX2 mux_inst_1330 (
  .O(mux_o_1330),
  .I0(mux_o_1058),
  .I1(mux_o_1059),
  .S0(ad[5])
);
MUX2 mux_inst_1331 (
  .O(mux_o_1331),
  .I0(mux_o_1060),
  .I1(mux_o_1061),
  .S0(ad[5])
);
MUX2 mux_inst_1332 (
  .O(mux_o_1332),
  .I0(mux_o_1062),
  .I1(mux_o_1063),
  .S0(ad[5])
);
MUX2 mux_inst_1333 (
  .O(mux_o_1333),
  .I0(mux_o_1064),
  .I1(mux_o_1065),
  .S0(ad[5])
);
MUX2 mux_inst_1334 (
  .O(mux_o_1334),
  .I0(mux_o_1066),
  .I1(mux_o_1067),
  .S0(ad[5])
);
MUX2 mux_inst_1335 (
  .O(mux_o_1335),
  .I0(mux_o_1068),
  .I1(mux_o_1069),
  .S0(ad[5])
);
MUX2 mux_inst_1336 (
  .O(mux_o_1336),
  .I0(mux_o_1070),
  .I1(mux_o_1071),
  .S0(ad[5])
);
MUX2 mux_inst_1337 (
  .O(mux_o_1337),
  .I0(mux_o_1072),
  .I1(mux_o_1073),
  .S0(ad[5])
);
MUX2 mux_inst_1338 (
  .O(mux_o_1338),
  .I0(mux_o_1074),
  .I1(mux_o_1075),
  .S0(ad[5])
);
MUX2 mux_inst_1339 (
  .O(mux_o_1339),
  .I0(mux_o_1076),
  .I1(mux_o_1077),
  .S0(ad[5])
);
MUX2 mux_inst_1340 (
  .O(mux_o_1340),
  .I0(mux_o_1078),
  .I1(mux_o_1079),
  .S0(ad[5])
);
MUX2 mux_inst_1341 (
  .O(mux_o_1341),
  .I0(mux_o_1080),
  .I1(mux_o_1081),
  .S0(ad[5])
);
MUX2 mux_inst_1342 (
  .O(mux_o_1342),
  .I0(mux_o_1082),
  .I1(mux_o_1083),
  .S0(ad[5])
);
MUX2 mux_inst_1343 (
  .O(mux_o_1343),
  .I0(mux_o_1084),
  .I1(mux_o_1085),
  .S0(ad[5])
);
MUX2 mux_inst_1344 (
  .O(mux_o_1344),
  .I0(mux_o_1086),
  .I1(mux_o_1087),
  .S0(ad[5])
);
MUX2 mux_inst_1345 (
  .O(mux_o_1345),
  .I0(mux_o_1088),
  .I1(mux_o_1089),
  .S0(ad[5])
);
MUX2 mux_inst_1346 (
  .O(mux_o_1346),
  .I0(mux_o_1090),
  .I1(mux_o_1091),
  .S0(ad[5])
);
MUX2 mux_inst_1347 (
  .O(mux_o_1347),
  .I0(mux_o_1092),
  .I1(mux_o_1093),
  .S0(ad[5])
);
MUX2 mux_inst_1348 (
  .O(mux_o_1348),
  .I0(mux_o_1094),
  .I1(mux_o_1095),
  .S0(ad[5])
);
MUX2 mux_inst_1349 (
  .O(mux_o_1349),
  .I0(mux_o_1096),
  .I1(mux_o_1097),
  .S0(ad[5])
);
MUX2 mux_inst_1350 (
  .O(mux_o_1350),
  .I0(mux_o_1098),
  .I1(mux_o_1099),
  .S0(ad[5])
);
MUX2 mux_inst_1351 (
  .O(mux_o_1351),
  .I0(mux_o_1100),
  .I1(mux_o_1101),
  .S0(ad[5])
);
MUX2 mux_inst_1352 (
  .O(mux_o_1352),
  .I0(mux_o_1102),
  .I1(mux_o_1103),
  .S0(ad[5])
);
MUX2 mux_inst_1353 (
  .O(mux_o_1353),
  .I0(mux_o_1104),
  .I1(mux_o_1105),
  .S0(ad[5])
);
MUX2 mux_inst_1354 (
  .O(mux_o_1354),
  .I0(mux_o_1106),
  .I1(mux_o_1107),
  .S0(ad[5])
);
MUX2 mux_inst_1355 (
  .O(mux_o_1355),
  .I0(mux_o_1108),
  .I1(mux_o_1109),
  .S0(ad[5])
);
MUX2 mux_inst_1356 (
  .O(mux_o_1356),
  .I0(mux_o_1110),
  .I1(mux_o_1111),
  .S0(ad[5])
);
MUX2 mux_inst_1357 (
  .O(mux_o_1357),
  .I0(mux_o_1112),
  .I1(mux_o_1113),
  .S0(ad[5])
);
MUX2 mux_inst_1358 (
  .O(mux_o_1358),
  .I0(mux_o_1114),
  .I1(mux_o_1115),
  .S0(ad[5])
);
MUX2 mux_inst_1359 (
  .O(mux_o_1359),
  .I0(mux_o_1116),
  .I1(mux_o_1117),
  .S0(ad[5])
);
MUX2 mux_inst_1360 (
  .O(mux_o_1360),
  .I0(mux_o_1118),
  .I1(mux_o_1119),
  .S0(ad[5])
);
MUX2 mux_inst_1361 (
  .O(mux_o_1361),
  .I0(mux_o_1120),
  .I1(mux_o_1121),
  .S0(ad[5])
);
MUX2 mux_inst_1362 (
  .O(mux_o_1362),
  .I0(mux_o_1122),
  .I1(mux_o_1123),
  .S0(ad[5])
);
MUX2 mux_inst_1363 (
  .O(mux_o_1363),
  .I0(mux_o_1124),
  .I1(mux_o_1125),
  .S0(ad[5])
);
MUX2 mux_inst_1364 (
  .O(mux_o_1364),
  .I0(mux_o_1126),
  .I1(mux_o_1127),
  .S0(ad[5])
);
MUX2 mux_inst_1365 (
  .O(mux_o_1365),
  .I0(mux_o_1128),
  .I1(mux_o_1129),
  .S0(ad[5])
);
MUX2 mux_inst_1366 (
  .O(mux_o_1366),
  .I0(mux_o_1130),
  .I1(mux_o_1131),
  .S0(ad[5])
);
MUX2 mux_inst_1367 (
  .O(mux_o_1367),
  .I0(mux_o_1132),
  .I1(mux_o_1133),
  .S0(ad[5])
);
MUX2 mux_inst_1368 (
  .O(mux_o_1368),
  .I0(mux_o_1134),
  .I1(mux_o_1135),
  .S0(ad[5])
);
MUX2 mux_inst_1369 (
  .O(mux_o_1369),
  .I0(mux_o_1136),
  .I1(mux_o_1137),
  .S0(ad[5])
);
MUX2 mux_inst_1370 (
  .O(mux_o_1370),
  .I0(mux_o_1138),
  .I1(mux_o_1139),
  .S0(ad[5])
);
MUX2 mux_inst_1371 (
  .O(mux_o_1371),
  .I0(mux_o_1140),
  .I1(mux_o_1141),
  .S0(ad[5])
);
MUX2 mux_inst_1372 (
  .O(mux_o_1372),
  .I0(mux_o_1142),
  .I1(mux_o_1143),
  .S0(ad[5])
);
MUX2 mux_inst_1373 (
  .O(mux_o_1373),
  .I0(mux_o_1144),
  .I1(mux_o_1145),
  .S0(ad[5])
);
MUX2 mux_inst_1374 (
  .O(mux_o_1374),
  .I0(mux_o_1146),
  .I1(mux_o_1147),
  .S0(ad[5])
);
MUX2 mux_inst_1375 (
  .O(mux_o_1375),
  .I0(mux_o_1148),
  .I1(mux_o_1149),
  .S0(ad[5])
);
MUX2 mux_inst_1376 (
  .O(mux_o_1376),
  .I0(mux_o_1150),
  .I1(mux_o_1151),
  .S0(ad[5])
);
MUX2 mux_inst_1377 (
  .O(mux_o_1377),
  .I0(mux_o_1152),
  .I1(mux_o_1153),
  .S0(ad[5])
);
MUX2 mux_inst_1378 (
  .O(mux_o_1378),
  .I0(mux_o_1154),
  .I1(mux_o_1155),
  .S0(ad[5])
);
MUX2 mux_inst_1379 (
  .O(mux_o_1379),
  .I0(mux_o_1156),
  .I1(mux_o_1157),
  .S0(ad[5])
);
MUX2 mux_inst_1380 (
  .O(mux_o_1380),
  .I0(mux_o_1158),
  .I1(mux_o_1159),
  .S0(ad[5])
);
MUX2 mux_inst_1381 (
  .O(mux_o_1381),
  .I0(mux_o_1160),
  .I1(mux_o_1161),
  .S0(ad[5])
);
MUX2 mux_inst_1382 (
  .O(mux_o_1382),
  .I0(mux_o_1162),
  .I1(mux_o_1163),
  .S0(ad[5])
);
MUX2 mux_inst_1383 (
  .O(mux_o_1383),
  .I0(mux_o_1164),
  .I1(mux_o_1165),
  .S0(ad[5])
);
MUX2 mux_inst_1384 (
  .O(mux_o_1384),
  .I0(mux_o_1166),
  .I1(mux_o_1167),
  .S0(ad[5])
);
MUX2 mux_inst_1385 (
  .O(mux_o_1385),
  .I0(mux_o_1168),
  .I1(mux_o_1169),
  .S0(ad[5])
);
MUX2 mux_inst_1386 (
  .O(mux_o_1386),
  .I0(mux_o_1170),
  .I1(mux_o_1171),
  .S0(ad[5])
);
MUX2 mux_inst_1387 (
  .O(mux_o_1387),
  .I0(mux_o_1172),
  .I1(mux_o_1173),
  .S0(ad[5])
);
MUX2 mux_inst_1388 (
  .O(mux_o_1388),
  .I0(mux_o_1174),
  .I1(mux_o_1175),
  .S0(ad[5])
);
MUX2 mux_inst_1389 (
  .O(mux_o_1389),
  .I0(mux_o_1176),
  .I1(mux_o_1177),
  .S0(ad[5])
);
MUX2 mux_inst_1390 (
  .O(mux_o_1390),
  .I0(mux_o_1178),
  .I1(mux_o_1179),
  .S0(ad[5])
);
MUX2 mux_inst_1391 (
  .O(mux_o_1391),
  .I0(mux_o_1180),
  .I1(mux_o_1181),
  .S0(ad[5])
);
MUX2 mux_inst_1392 (
  .O(mux_o_1392),
  .I0(mux_o_1182),
  .I1(mux_o_1183),
  .S0(ad[5])
);
MUX2 mux_inst_1393 (
  .O(mux_o_1393),
  .I0(mux_o_1184),
  .I1(mux_o_1185),
  .S0(ad[5])
);
MUX2 mux_inst_1394 (
  .O(mux_o_1394),
  .I0(mux_o_1186),
  .I1(mux_o_1187),
  .S0(ad[5])
);
MUX2 mux_inst_1395 (
  .O(mux_o_1395),
  .I0(mux_o_1188),
  .I1(mux_o_1189),
  .S0(ad[5])
);
MUX2 mux_inst_1396 (
  .O(mux_o_1396),
  .I0(mux_o_1190),
  .I1(mux_o_1191),
  .S0(ad[5])
);
MUX2 mux_inst_1397 (
  .O(mux_o_1397),
  .I0(mux_o_1192),
  .I1(mux_o_1193),
  .S0(ad[5])
);
MUX2 mux_inst_1398 (
  .O(mux_o_1398),
  .I0(mux_o_1194),
  .I1(mux_o_1195),
  .S0(ad[5])
);
MUX2 mux_inst_1399 (
  .O(mux_o_1399),
  .I0(mux_o_1196),
  .I1(mux_o_1197),
  .S0(ad[5])
);
MUX2 mux_inst_1400 (
  .O(mux_o_1400),
  .I0(mux_o_1198),
  .I1(mux_o_1199),
  .S0(ad[5])
);
MUX2 mux_inst_1401 (
  .O(mux_o_1401),
  .I0(mux_o_1200),
  .I1(mux_o_1201),
  .S0(ad[5])
);
MUX2 mux_inst_1402 (
  .O(mux_o_1402),
  .I0(mux_o_1202),
  .I1(mux_o_1203),
  .S0(ad[6])
);
MUX2 mux_inst_1403 (
  .O(mux_o_1403),
  .I0(mux_o_1204),
  .I1(mux_o_1205),
  .S0(ad[6])
);
MUX2 mux_inst_1404 (
  .O(mux_o_1404),
  .I0(mux_o_1206),
  .I1(mux_o_1207),
  .S0(ad[6])
);
MUX2 mux_inst_1405 (
  .O(mux_o_1405),
  .I0(mux_o_1208),
  .I1(mux_o_1209),
  .S0(ad[6])
);
MUX2 mux_inst_1406 (
  .O(mux_o_1406),
  .I0(mux_o_1210),
  .I1(mux_o_1211),
  .S0(ad[6])
);
MUX2 mux_inst_1407 (
  .O(mux_o_1407),
  .I0(mux_o_1212),
  .I1(mux_o_1213),
  .S0(ad[6])
);
MUX2 mux_inst_1408 (
  .O(mux_o_1408),
  .I0(mux_o_1214),
  .I1(mux_o_1215),
  .S0(ad[6])
);
MUX2 mux_inst_1409 (
  .O(mux_o_1409),
  .I0(mux_o_1216),
  .I1(mux_o_1217),
  .S0(ad[6])
);
MUX2 mux_inst_1410 (
  .O(mux_o_1410),
  .I0(mux_o_1218),
  .I1(mux_o_1219),
  .S0(ad[6])
);
MUX2 mux_inst_1411 (
  .O(mux_o_1411),
  .I0(mux_o_1220),
  .I1(mux_o_1221),
  .S0(ad[6])
);
MUX2 mux_inst_1412 (
  .O(mux_o_1412),
  .I0(mux_o_1222),
  .I1(mux_o_1223),
  .S0(ad[6])
);
MUX2 mux_inst_1413 (
  .O(mux_o_1413),
  .I0(mux_o_1224),
  .I1(mux_o_1225),
  .S0(ad[6])
);
MUX2 mux_inst_1414 (
  .O(mux_o_1414),
  .I0(mux_o_1226),
  .I1(mux_o_1227),
  .S0(ad[6])
);
MUX2 mux_inst_1415 (
  .O(mux_o_1415),
  .I0(mux_o_1228),
  .I1(mux_o_1229),
  .S0(ad[6])
);
MUX2 mux_inst_1416 (
  .O(mux_o_1416),
  .I0(mux_o_1230),
  .I1(mux_o_1231),
  .S0(ad[6])
);
MUX2 mux_inst_1417 (
  .O(mux_o_1417),
  .I0(mux_o_1232),
  .I1(mux_o_1233),
  .S0(ad[6])
);
MUX2 mux_inst_1418 (
  .O(mux_o_1418),
  .I0(mux_o_1234),
  .I1(mux_o_1235),
  .S0(ad[6])
);
MUX2 mux_inst_1419 (
  .O(mux_o_1419),
  .I0(mux_o_1236),
  .I1(mux_o_1237),
  .S0(ad[6])
);
MUX2 mux_inst_1420 (
  .O(mux_o_1420),
  .I0(mux_o_1238),
  .I1(mux_o_1239),
  .S0(ad[6])
);
MUX2 mux_inst_1421 (
  .O(mux_o_1421),
  .I0(mux_o_1240),
  .I1(mux_o_1241),
  .S0(ad[6])
);
MUX2 mux_inst_1422 (
  .O(mux_o_1422),
  .I0(mux_o_1242),
  .I1(mux_o_1243),
  .S0(ad[6])
);
MUX2 mux_inst_1423 (
  .O(mux_o_1423),
  .I0(mux_o_1244),
  .I1(mux_o_1245),
  .S0(ad[6])
);
MUX2 mux_inst_1424 (
  .O(mux_o_1424),
  .I0(mux_o_1246),
  .I1(mux_o_1247),
  .S0(ad[6])
);
MUX2 mux_inst_1425 (
  .O(mux_o_1425),
  .I0(mux_o_1248),
  .I1(mux_o_1249),
  .S0(ad[6])
);
MUX2 mux_inst_1426 (
  .O(mux_o_1426),
  .I0(mux_o_1250),
  .I1(mux_o_1251),
  .S0(ad[6])
);
MUX2 mux_inst_1427 (
  .O(mux_o_1427),
  .I0(mux_o_1252),
  .I1(mux_o_1253),
  .S0(ad[6])
);
MUX2 mux_inst_1428 (
  .O(mux_o_1428),
  .I0(mux_o_1254),
  .I1(mux_o_1255),
  .S0(ad[6])
);
MUX2 mux_inst_1429 (
  .O(mux_o_1429),
  .I0(mux_o_1256),
  .I1(mux_o_1257),
  .S0(ad[6])
);
MUX2 mux_inst_1430 (
  .O(mux_o_1430),
  .I0(mux_o_1258),
  .I1(mux_o_1259),
  .S0(ad[6])
);
MUX2 mux_inst_1431 (
  .O(mux_o_1431),
  .I0(mux_o_1260),
  .I1(mux_o_1261),
  .S0(ad[6])
);
MUX2 mux_inst_1432 (
  .O(mux_o_1432),
  .I0(mux_o_1262),
  .I1(mux_o_1263),
  .S0(ad[6])
);
MUX2 mux_inst_1433 (
  .O(mux_o_1433),
  .I0(mux_o_1264),
  .I1(mux_o_1265),
  .S0(ad[6])
);
MUX2 mux_inst_1434 (
  .O(mux_o_1434),
  .I0(mux_o_1266),
  .I1(mux_o_1267),
  .S0(ad[6])
);
MUX2 mux_inst_1435 (
  .O(mux_o_1435),
  .I0(mux_o_1268),
  .I1(mux_o_1269),
  .S0(ad[6])
);
MUX2 mux_inst_1436 (
  .O(mux_o_1436),
  .I0(mux_o_1270),
  .I1(mux_o_1271),
  .S0(ad[6])
);
MUX2 mux_inst_1437 (
  .O(mux_o_1437),
  .I0(mux_o_1272),
  .I1(mux_o_1273),
  .S0(ad[6])
);
MUX2 mux_inst_1438 (
  .O(mux_o_1438),
  .I0(mux_o_1274),
  .I1(mux_o_1275),
  .S0(ad[6])
);
MUX2 mux_inst_1439 (
  .O(mux_o_1439),
  .I0(mux_o_1276),
  .I1(mux_o_1277),
  .S0(ad[6])
);
MUX2 mux_inst_1440 (
  .O(mux_o_1440),
  .I0(mux_o_1278),
  .I1(mux_o_1279),
  .S0(ad[6])
);
MUX2 mux_inst_1441 (
  .O(mux_o_1441),
  .I0(mux_o_1280),
  .I1(mux_o_1281),
  .S0(ad[6])
);
MUX2 mux_inst_1442 (
  .O(mux_o_1442),
  .I0(mux_o_1282),
  .I1(mux_o_1283),
  .S0(ad[6])
);
MUX2 mux_inst_1443 (
  .O(mux_o_1443),
  .I0(mux_o_1284),
  .I1(mux_o_1285),
  .S0(ad[6])
);
MUX2 mux_inst_1444 (
  .O(mux_o_1444),
  .I0(mux_o_1286),
  .I1(mux_o_1287),
  .S0(ad[6])
);
MUX2 mux_inst_1445 (
  .O(mux_o_1445),
  .I0(mux_o_1288),
  .I1(mux_o_1289),
  .S0(ad[6])
);
MUX2 mux_inst_1446 (
  .O(mux_o_1446),
  .I0(mux_o_1290),
  .I1(mux_o_1291),
  .S0(ad[6])
);
MUX2 mux_inst_1447 (
  .O(mux_o_1447),
  .I0(mux_o_1292),
  .I1(mux_o_1293),
  .S0(ad[6])
);
MUX2 mux_inst_1448 (
  .O(mux_o_1448),
  .I0(mux_o_1294),
  .I1(mux_o_1295),
  .S0(ad[6])
);
MUX2 mux_inst_1449 (
  .O(mux_o_1449),
  .I0(mux_o_1296),
  .I1(mux_o_1297),
  .S0(ad[6])
);
MUX2 mux_inst_1450 (
  .O(mux_o_1450),
  .I0(mux_o_1298),
  .I1(mux_o_1299),
  .S0(ad[6])
);
MUX2 mux_inst_1451 (
  .O(mux_o_1451),
  .I0(mux_o_1300),
  .I1(mux_o_1301),
  .S0(ad[6])
);
MUX2 mux_inst_1452 (
  .O(mux_o_1452),
  .I0(mux_o_1302),
  .I1(mux_o_1303),
  .S0(ad[6])
);
MUX2 mux_inst_1453 (
  .O(mux_o_1453),
  .I0(mux_o_1304),
  .I1(mux_o_1305),
  .S0(ad[6])
);
MUX2 mux_inst_1454 (
  .O(mux_o_1454),
  .I0(mux_o_1306),
  .I1(mux_o_1307),
  .S0(ad[6])
);
MUX2 mux_inst_1455 (
  .O(mux_o_1455),
  .I0(mux_o_1308),
  .I1(mux_o_1309),
  .S0(ad[6])
);
MUX2 mux_inst_1456 (
  .O(mux_o_1456),
  .I0(mux_o_1310),
  .I1(mux_o_1311),
  .S0(ad[6])
);
MUX2 mux_inst_1457 (
  .O(mux_o_1457),
  .I0(mux_o_1312),
  .I1(mux_o_1313),
  .S0(ad[6])
);
MUX2 mux_inst_1458 (
  .O(mux_o_1458),
  .I0(mux_o_1314),
  .I1(mux_o_1315),
  .S0(ad[6])
);
MUX2 mux_inst_1459 (
  .O(mux_o_1459),
  .I0(mux_o_1316),
  .I1(mux_o_1317),
  .S0(ad[6])
);
MUX2 mux_inst_1460 (
  .O(mux_o_1460),
  .I0(mux_o_1318),
  .I1(mux_o_1319),
  .S0(ad[6])
);
MUX2 mux_inst_1461 (
  .O(mux_o_1461),
  .I0(mux_o_1320),
  .I1(mux_o_1321),
  .S0(ad[6])
);
MUX2 mux_inst_1462 (
  .O(mux_o_1462),
  .I0(mux_o_1322),
  .I1(mux_o_1323),
  .S0(ad[6])
);
MUX2 mux_inst_1463 (
  .O(mux_o_1463),
  .I0(mux_o_1324),
  .I1(mux_o_1325),
  .S0(ad[6])
);
MUX2 mux_inst_1464 (
  .O(mux_o_1464),
  .I0(mux_o_1326),
  .I1(mux_o_1327),
  .S0(ad[6])
);
MUX2 mux_inst_1465 (
  .O(mux_o_1465),
  .I0(mux_o_1328),
  .I1(mux_o_1329),
  .S0(ad[6])
);
MUX2 mux_inst_1466 (
  .O(mux_o_1466),
  .I0(mux_o_1330),
  .I1(mux_o_1331),
  .S0(ad[6])
);
MUX2 mux_inst_1467 (
  .O(mux_o_1467),
  .I0(mux_o_1332),
  .I1(mux_o_1333),
  .S0(ad[6])
);
MUX2 mux_inst_1468 (
  .O(mux_o_1468),
  .I0(mux_o_1334),
  .I1(mux_o_1335),
  .S0(ad[6])
);
MUX2 mux_inst_1469 (
  .O(mux_o_1469),
  .I0(mux_o_1336),
  .I1(mux_o_1337),
  .S0(ad[6])
);
MUX2 mux_inst_1470 (
  .O(mux_o_1470),
  .I0(mux_o_1338),
  .I1(mux_o_1339),
  .S0(ad[6])
);
MUX2 mux_inst_1471 (
  .O(mux_o_1471),
  .I0(mux_o_1340),
  .I1(mux_o_1341),
  .S0(ad[6])
);
MUX2 mux_inst_1472 (
  .O(mux_o_1472),
  .I0(mux_o_1342),
  .I1(mux_o_1343),
  .S0(ad[6])
);
MUX2 mux_inst_1473 (
  .O(mux_o_1473),
  .I0(mux_o_1344),
  .I1(mux_o_1345),
  .S0(ad[6])
);
MUX2 mux_inst_1474 (
  .O(mux_o_1474),
  .I0(mux_o_1346),
  .I1(mux_o_1347),
  .S0(ad[6])
);
MUX2 mux_inst_1475 (
  .O(mux_o_1475),
  .I0(mux_o_1348),
  .I1(mux_o_1349),
  .S0(ad[6])
);
MUX2 mux_inst_1476 (
  .O(mux_o_1476),
  .I0(mux_o_1350),
  .I1(mux_o_1351),
  .S0(ad[6])
);
MUX2 mux_inst_1477 (
  .O(mux_o_1477),
  .I0(mux_o_1352),
  .I1(mux_o_1353),
  .S0(ad[6])
);
MUX2 mux_inst_1478 (
  .O(mux_o_1478),
  .I0(mux_o_1354),
  .I1(mux_o_1355),
  .S0(ad[6])
);
MUX2 mux_inst_1479 (
  .O(mux_o_1479),
  .I0(mux_o_1356),
  .I1(mux_o_1357),
  .S0(ad[6])
);
MUX2 mux_inst_1480 (
  .O(mux_o_1480),
  .I0(mux_o_1358),
  .I1(mux_o_1359),
  .S0(ad[6])
);
MUX2 mux_inst_1481 (
  .O(mux_o_1481),
  .I0(mux_o_1360),
  .I1(mux_o_1361),
  .S0(ad[6])
);
MUX2 mux_inst_1482 (
  .O(mux_o_1482),
  .I0(mux_o_1362),
  .I1(mux_o_1363),
  .S0(ad[6])
);
MUX2 mux_inst_1483 (
  .O(mux_o_1483),
  .I0(mux_o_1364),
  .I1(mux_o_1365),
  .S0(ad[6])
);
MUX2 mux_inst_1484 (
  .O(mux_o_1484),
  .I0(mux_o_1366),
  .I1(mux_o_1367),
  .S0(ad[6])
);
MUX2 mux_inst_1485 (
  .O(mux_o_1485),
  .I0(mux_o_1368),
  .I1(mux_o_1369),
  .S0(ad[6])
);
MUX2 mux_inst_1486 (
  .O(mux_o_1486),
  .I0(mux_o_1370),
  .I1(mux_o_1371),
  .S0(ad[6])
);
MUX2 mux_inst_1487 (
  .O(mux_o_1487),
  .I0(mux_o_1372),
  .I1(mux_o_1373),
  .S0(ad[6])
);
MUX2 mux_inst_1488 (
  .O(mux_o_1488),
  .I0(mux_o_1374),
  .I1(mux_o_1375),
  .S0(ad[6])
);
MUX2 mux_inst_1489 (
  .O(mux_o_1489),
  .I0(mux_o_1376),
  .I1(mux_o_1377),
  .S0(ad[6])
);
MUX2 mux_inst_1490 (
  .O(mux_o_1490),
  .I0(mux_o_1378),
  .I1(mux_o_1379),
  .S0(ad[6])
);
MUX2 mux_inst_1491 (
  .O(mux_o_1491),
  .I0(mux_o_1380),
  .I1(mux_o_1381),
  .S0(ad[6])
);
MUX2 mux_inst_1492 (
  .O(mux_o_1492),
  .I0(mux_o_1382),
  .I1(mux_o_1383),
  .S0(ad[6])
);
MUX2 mux_inst_1493 (
  .O(mux_o_1493),
  .I0(mux_o_1384),
  .I1(mux_o_1385),
  .S0(ad[6])
);
MUX2 mux_inst_1494 (
  .O(mux_o_1494),
  .I0(mux_o_1386),
  .I1(mux_o_1387),
  .S0(ad[6])
);
MUX2 mux_inst_1495 (
  .O(mux_o_1495),
  .I0(mux_o_1388),
  .I1(mux_o_1389),
  .S0(ad[6])
);
MUX2 mux_inst_1496 (
  .O(mux_o_1496),
  .I0(mux_o_1390),
  .I1(mux_o_1391),
  .S0(ad[6])
);
MUX2 mux_inst_1497 (
  .O(mux_o_1497),
  .I0(mux_o_1392),
  .I1(mux_o_1393),
  .S0(ad[6])
);
MUX2 mux_inst_1498 (
  .O(mux_o_1498),
  .I0(mux_o_1394),
  .I1(mux_o_1395),
  .S0(ad[6])
);
MUX2 mux_inst_1499 (
  .O(mux_o_1499),
  .I0(mux_o_1396),
  .I1(mux_o_1397),
  .S0(ad[6])
);
MUX2 mux_inst_1500 (
  .O(mux_o_1500),
  .I0(mux_o_1398),
  .I1(mux_o_1399),
  .S0(ad[6])
);
MUX2 mux_inst_1501 (
  .O(mux_o_1501),
  .I0(mux_o_1400),
  .I1(mux_o_1401),
  .S0(ad[6])
);
MUX2 mux_inst_1502 (
  .O(mux_o_1502),
  .I0(mux_o_1402),
  .I1(mux_o_1403),
  .S0(ad[7])
);
MUX2 mux_inst_1503 (
  .O(mux_o_1503),
  .I0(mux_o_1404),
  .I1(mux_o_1405),
  .S0(ad[7])
);
MUX2 mux_inst_1504 (
  .O(mux_o_1504),
  .I0(mux_o_1406),
  .I1(mux_o_1407),
  .S0(ad[7])
);
MUX2 mux_inst_1505 (
  .O(mux_o_1505),
  .I0(mux_o_1408),
  .I1(mux_o_1409),
  .S0(ad[7])
);
MUX2 mux_inst_1506 (
  .O(mux_o_1506),
  .I0(mux_o_1410),
  .I1(mux_o_1411),
  .S0(ad[7])
);
MUX2 mux_inst_1507 (
  .O(mux_o_1507),
  .I0(mux_o_1412),
  .I1(mux_o_1413),
  .S0(ad[7])
);
MUX2 mux_inst_1508 (
  .O(mux_o_1508),
  .I0(mux_o_1414),
  .I1(mux_o_1415),
  .S0(ad[7])
);
MUX2 mux_inst_1509 (
  .O(mux_o_1509),
  .I0(mux_o_1416),
  .I1(mux_o_1417),
  .S0(ad[7])
);
MUX2 mux_inst_1510 (
  .O(mux_o_1510),
  .I0(mux_o_1418),
  .I1(mux_o_1419),
  .S0(ad[7])
);
MUX2 mux_inst_1511 (
  .O(mux_o_1511),
  .I0(mux_o_1420),
  .I1(mux_o_1421),
  .S0(ad[7])
);
MUX2 mux_inst_1512 (
  .O(mux_o_1512),
  .I0(mux_o_1422),
  .I1(mux_o_1423),
  .S0(ad[7])
);
MUX2 mux_inst_1513 (
  .O(mux_o_1513),
  .I0(mux_o_1424),
  .I1(mux_o_1425),
  .S0(ad[7])
);
MUX2 mux_inst_1514 (
  .O(mux_o_1514),
  .I0(mux_o_1426),
  .I1(mux_o_1427),
  .S0(ad[7])
);
MUX2 mux_inst_1515 (
  .O(mux_o_1515),
  .I0(mux_o_1428),
  .I1(mux_o_1429),
  .S0(ad[7])
);
MUX2 mux_inst_1516 (
  .O(mux_o_1516),
  .I0(mux_o_1430),
  .I1(mux_o_1431),
  .S0(ad[7])
);
MUX2 mux_inst_1517 (
  .O(mux_o_1517),
  .I0(mux_o_1432),
  .I1(mux_o_1433),
  .S0(ad[7])
);
MUX2 mux_inst_1518 (
  .O(mux_o_1518),
  .I0(mux_o_1434),
  .I1(mux_o_1435),
  .S0(ad[7])
);
MUX2 mux_inst_1519 (
  .O(mux_o_1519),
  .I0(mux_o_1436),
  .I1(mux_o_1437),
  .S0(ad[7])
);
MUX2 mux_inst_1520 (
  .O(mux_o_1520),
  .I0(mux_o_1438),
  .I1(mux_o_1439),
  .S0(ad[7])
);
MUX2 mux_inst_1521 (
  .O(mux_o_1521),
  .I0(mux_o_1440),
  .I1(mux_o_1441),
  .S0(ad[7])
);
MUX2 mux_inst_1522 (
  .O(mux_o_1522),
  .I0(mux_o_1442),
  .I1(mux_o_1443),
  .S0(ad[7])
);
MUX2 mux_inst_1523 (
  .O(mux_o_1523),
  .I0(mux_o_1444),
  .I1(mux_o_1445),
  .S0(ad[7])
);
MUX2 mux_inst_1524 (
  .O(mux_o_1524),
  .I0(mux_o_1446),
  .I1(mux_o_1447),
  .S0(ad[7])
);
MUX2 mux_inst_1525 (
  .O(mux_o_1525),
  .I0(mux_o_1448),
  .I1(mux_o_1449),
  .S0(ad[7])
);
MUX2 mux_inst_1526 (
  .O(mux_o_1526),
  .I0(mux_o_1450),
  .I1(mux_o_1451),
  .S0(ad[7])
);
MUX2 mux_inst_1527 (
  .O(mux_o_1527),
  .I0(mux_o_1452),
  .I1(mux_o_1453),
  .S0(ad[7])
);
MUX2 mux_inst_1528 (
  .O(mux_o_1528),
  .I0(mux_o_1454),
  .I1(mux_o_1455),
  .S0(ad[7])
);
MUX2 mux_inst_1529 (
  .O(mux_o_1529),
  .I0(mux_o_1456),
  .I1(mux_o_1457),
  .S0(ad[7])
);
MUX2 mux_inst_1530 (
  .O(mux_o_1530),
  .I0(mux_o_1458),
  .I1(mux_o_1459),
  .S0(ad[7])
);
MUX2 mux_inst_1531 (
  .O(mux_o_1531),
  .I0(mux_o_1460),
  .I1(mux_o_1461),
  .S0(ad[7])
);
MUX2 mux_inst_1532 (
  .O(mux_o_1532),
  .I0(mux_o_1462),
  .I1(mux_o_1463),
  .S0(ad[7])
);
MUX2 mux_inst_1533 (
  .O(mux_o_1533),
  .I0(mux_o_1464),
  .I1(mux_o_1465),
  .S0(ad[7])
);
MUX2 mux_inst_1534 (
  .O(mux_o_1534),
  .I0(mux_o_1466),
  .I1(mux_o_1467),
  .S0(ad[7])
);
MUX2 mux_inst_1535 (
  .O(mux_o_1535),
  .I0(mux_o_1468),
  .I1(mux_o_1469),
  .S0(ad[7])
);
MUX2 mux_inst_1536 (
  .O(mux_o_1536),
  .I0(mux_o_1470),
  .I1(mux_o_1471),
  .S0(ad[7])
);
MUX2 mux_inst_1537 (
  .O(mux_o_1537),
  .I0(mux_o_1472),
  .I1(mux_o_1473),
  .S0(ad[7])
);
MUX2 mux_inst_1538 (
  .O(mux_o_1538),
  .I0(mux_o_1474),
  .I1(mux_o_1475),
  .S0(ad[7])
);
MUX2 mux_inst_1539 (
  .O(mux_o_1539),
  .I0(mux_o_1476),
  .I1(mux_o_1477),
  .S0(ad[7])
);
MUX2 mux_inst_1540 (
  .O(mux_o_1540),
  .I0(mux_o_1478),
  .I1(mux_o_1479),
  .S0(ad[7])
);
MUX2 mux_inst_1541 (
  .O(mux_o_1541),
  .I0(mux_o_1480),
  .I1(mux_o_1481),
  .S0(ad[7])
);
MUX2 mux_inst_1542 (
  .O(mux_o_1542),
  .I0(mux_o_1482),
  .I1(mux_o_1483),
  .S0(ad[7])
);
MUX2 mux_inst_1543 (
  .O(mux_o_1543),
  .I0(mux_o_1484),
  .I1(mux_o_1485),
  .S0(ad[7])
);
MUX2 mux_inst_1544 (
  .O(mux_o_1544),
  .I0(mux_o_1486),
  .I1(mux_o_1487),
  .S0(ad[7])
);
MUX2 mux_inst_1545 (
  .O(mux_o_1545),
  .I0(mux_o_1488),
  .I1(mux_o_1489),
  .S0(ad[7])
);
MUX2 mux_inst_1546 (
  .O(mux_o_1546),
  .I0(mux_o_1490),
  .I1(mux_o_1491),
  .S0(ad[7])
);
MUX2 mux_inst_1547 (
  .O(mux_o_1547),
  .I0(mux_o_1492),
  .I1(mux_o_1493),
  .S0(ad[7])
);
MUX2 mux_inst_1548 (
  .O(mux_o_1548),
  .I0(mux_o_1494),
  .I1(mux_o_1495),
  .S0(ad[7])
);
MUX2 mux_inst_1549 (
  .O(mux_o_1549),
  .I0(mux_o_1496),
  .I1(mux_o_1497),
  .S0(ad[7])
);
MUX2 mux_inst_1550 (
  .O(mux_o_1550),
  .I0(mux_o_1498),
  .I1(mux_o_1499),
  .S0(ad[7])
);
MUX2 mux_inst_1551 (
  .O(mux_o_1551),
  .I0(mux_o_1500),
  .I1(mux_o_1501),
  .S0(ad[7])
);
MUX2 mux_inst_1552 (
  .O(mux_o_1552),
  .I0(mux_o_1502),
  .I1(mux_o_1503),
  .S0(ad[8])
);
MUX2 mux_inst_1553 (
  .O(mux_o_1553),
  .I0(mux_o_1504),
  .I1(mux_o_1505),
  .S0(ad[8])
);
MUX2 mux_inst_1554 (
  .O(mux_o_1554),
  .I0(mux_o_1506),
  .I1(mux_o_1507),
  .S0(ad[8])
);
MUX2 mux_inst_1555 (
  .O(mux_o_1555),
  .I0(mux_o_1508),
  .I1(mux_o_1509),
  .S0(ad[8])
);
MUX2 mux_inst_1556 (
  .O(mux_o_1556),
  .I0(mux_o_1510),
  .I1(mux_o_1511),
  .S0(ad[8])
);
MUX2 mux_inst_1557 (
  .O(mux_o_1557),
  .I0(mux_o_1512),
  .I1(mux_o_1513),
  .S0(ad[8])
);
MUX2 mux_inst_1558 (
  .O(mux_o_1558),
  .I0(mux_o_1514),
  .I1(mux_o_1515),
  .S0(ad[8])
);
MUX2 mux_inst_1559 (
  .O(mux_o_1559),
  .I0(mux_o_1516),
  .I1(mux_o_1517),
  .S0(ad[8])
);
MUX2 mux_inst_1560 (
  .O(mux_o_1560),
  .I0(mux_o_1518),
  .I1(mux_o_1519),
  .S0(ad[8])
);
MUX2 mux_inst_1561 (
  .O(mux_o_1561),
  .I0(mux_o_1520),
  .I1(mux_o_1521),
  .S0(ad[8])
);
MUX2 mux_inst_1562 (
  .O(mux_o_1562),
  .I0(mux_o_1522),
  .I1(mux_o_1523),
  .S0(ad[8])
);
MUX2 mux_inst_1563 (
  .O(mux_o_1563),
  .I0(mux_o_1524),
  .I1(mux_o_1525),
  .S0(ad[8])
);
MUX2 mux_inst_1564 (
  .O(mux_o_1564),
  .I0(mux_o_1526),
  .I1(mux_o_1527),
  .S0(ad[8])
);
MUX2 mux_inst_1565 (
  .O(mux_o_1565),
  .I0(mux_o_1528),
  .I1(mux_o_1529),
  .S0(ad[8])
);
MUX2 mux_inst_1566 (
  .O(mux_o_1566),
  .I0(mux_o_1530),
  .I1(mux_o_1531),
  .S0(ad[8])
);
MUX2 mux_inst_1567 (
  .O(mux_o_1567),
  .I0(mux_o_1532),
  .I1(mux_o_1533),
  .S0(ad[8])
);
MUX2 mux_inst_1568 (
  .O(mux_o_1568),
  .I0(mux_o_1534),
  .I1(mux_o_1535),
  .S0(ad[8])
);
MUX2 mux_inst_1569 (
  .O(mux_o_1569),
  .I0(mux_o_1536),
  .I1(mux_o_1537),
  .S0(ad[8])
);
MUX2 mux_inst_1570 (
  .O(mux_o_1570),
  .I0(mux_o_1538),
  .I1(mux_o_1539),
  .S0(ad[8])
);
MUX2 mux_inst_1571 (
  .O(mux_o_1571),
  .I0(mux_o_1540),
  .I1(mux_o_1541),
  .S0(ad[8])
);
MUX2 mux_inst_1572 (
  .O(mux_o_1572),
  .I0(mux_o_1542),
  .I1(mux_o_1543),
  .S0(ad[8])
);
MUX2 mux_inst_1573 (
  .O(mux_o_1573),
  .I0(mux_o_1544),
  .I1(mux_o_1545),
  .S0(ad[8])
);
MUX2 mux_inst_1574 (
  .O(mux_o_1574),
  .I0(mux_o_1546),
  .I1(mux_o_1547),
  .S0(ad[8])
);
MUX2 mux_inst_1575 (
  .O(mux_o_1575),
  .I0(mux_o_1548),
  .I1(mux_o_1549),
  .S0(ad[8])
);
MUX2 mux_inst_1576 (
  .O(mux_o_1576),
  .I0(mux_o_1550),
  .I1(mux_o_1551),
  .S0(ad[8])
);
MUX2 mux_inst_1577 (
  .O(mux_o_1577),
  .I0(mux_o_1552),
  .I1(mux_o_1553),
  .S0(ad[9])
);
MUX2 mux_inst_1578 (
  .O(mux_o_1578),
  .I0(mux_o_1554),
  .I1(mux_o_1555),
  .S0(ad[9])
);
MUX2 mux_inst_1579 (
  .O(mux_o_1579),
  .I0(mux_o_1556),
  .I1(mux_o_1557),
  .S0(ad[9])
);
MUX2 mux_inst_1580 (
  .O(mux_o_1580),
  .I0(mux_o_1558),
  .I1(mux_o_1559),
  .S0(ad[9])
);
MUX2 mux_inst_1581 (
  .O(mux_o_1581),
  .I0(mux_o_1560),
  .I1(mux_o_1561),
  .S0(ad[9])
);
MUX2 mux_inst_1582 (
  .O(mux_o_1582),
  .I0(mux_o_1562),
  .I1(mux_o_1563),
  .S0(ad[9])
);
MUX2 mux_inst_1583 (
  .O(mux_o_1583),
  .I0(mux_o_1564),
  .I1(mux_o_1565),
  .S0(ad[9])
);
MUX2 mux_inst_1584 (
  .O(mux_o_1584),
  .I0(mux_o_1566),
  .I1(mux_o_1567),
  .S0(ad[9])
);
MUX2 mux_inst_1585 (
  .O(mux_o_1585),
  .I0(mux_o_1568),
  .I1(mux_o_1569),
  .S0(ad[9])
);
MUX2 mux_inst_1586 (
  .O(mux_o_1586),
  .I0(mux_o_1570),
  .I1(mux_o_1571),
  .S0(ad[9])
);
MUX2 mux_inst_1587 (
  .O(mux_o_1587),
  .I0(mux_o_1572),
  .I1(mux_o_1573),
  .S0(ad[9])
);
MUX2 mux_inst_1588 (
  .O(mux_o_1588),
  .I0(mux_o_1574),
  .I1(mux_o_1575),
  .S0(ad[9])
);
MUX2 mux_inst_1590 (
  .O(mux_o_1590),
  .I0(mux_o_1577),
  .I1(mux_o_1578),
  .S0(ad[10])
);
MUX2 mux_inst_1591 (
  .O(mux_o_1591),
  .I0(mux_o_1579),
  .I1(mux_o_1580),
  .S0(ad[10])
);
MUX2 mux_inst_1592 (
  .O(mux_o_1592),
  .I0(mux_o_1581),
  .I1(mux_o_1582),
  .S0(ad[10])
);
MUX2 mux_inst_1593 (
  .O(mux_o_1593),
  .I0(mux_o_1583),
  .I1(mux_o_1584),
  .S0(ad[10])
);
MUX2 mux_inst_1594 (
  .O(mux_o_1594),
  .I0(mux_o_1585),
  .I1(mux_o_1586),
  .S0(ad[10])
);
MUX2 mux_inst_1595 (
  .O(mux_o_1595),
  .I0(mux_o_1587),
  .I1(mux_o_1588),
  .S0(ad[10])
);
MUX2 mux_inst_1597 (
  .O(mux_o_1597),
  .I0(mux_o_1590),
  .I1(mux_o_1591),
  .S0(ad[11])
);
MUX2 mux_inst_1598 (
  .O(mux_o_1598),
  .I0(mux_o_1592),
  .I1(mux_o_1593),
  .S0(ad[11])
);
MUX2 mux_inst_1599 (
  .O(mux_o_1599),
  .I0(mux_o_1594),
  .I1(mux_o_1595),
  .S0(ad[11])
);
MUX2 mux_inst_1601 (
  .O(mux_o_1601),
  .I0(mux_o_1597),
  .I1(mux_o_1598),
  .S0(ad[12])
);
MUX2 mux_inst_1602 (
  .O(mux_o_1602),
  .I0(mux_o_1599),
  .I1(mux_o_1576),
  .S0(ad[12])
);
MUX2 mux_inst_1603 (
  .O(dout[1]),
  .I0(mux_o_1601),
  .I1(mux_o_1602),
  .S0(ad[13])
);
MUX2 mux_inst_1604 (
  .O(mux_o_1604),
  .I0(ram16s_inst_0_dout[2]),
  .I1(ram16s_inst_1_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1605 (
  .O(mux_o_1605),
  .I0(ram16s_inst_2_dout[2]),
  .I1(ram16s_inst_3_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1606 (
  .O(mux_o_1606),
  .I0(ram16s_inst_4_dout[2]),
  .I1(ram16s_inst_5_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1607 (
  .O(mux_o_1607),
  .I0(ram16s_inst_6_dout[2]),
  .I1(ram16s_inst_7_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1608 (
  .O(mux_o_1608),
  .I0(ram16s_inst_8_dout[2]),
  .I1(ram16s_inst_9_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1609 (
  .O(mux_o_1609),
  .I0(ram16s_inst_10_dout[2]),
  .I1(ram16s_inst_11_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1610 (
  .O(mux_o_1610),
  .I0(ram16s_inst_12_dout[2]),
  .I1(ram16s_inst_13_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1611 (
  .O(mux_o_1611),
  .I0(ram16s_inst_14_dout[2]),
  .I1(ram16s_inst_15_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1612 (
  .O(mux_o_1612),
  .I0(ram16s_inst_16_dout[2]),
  .I1(ram16s_inst_17_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1613 (
  .O(mux_o_1613),
  .I0(ram16s_inst_18_dout[2]),
  .I1(ram16s_inst_19_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1614 (
  .O(mux_o_1614),
  .I0(ram16s_inst_20_dout[2]),
  .I1(ram16s_inst_21_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1615 (
  .O(mux_o_1615),
  .I0(ram16s_inst_22_dout[2]),
  .I1(ram16s_inst_23_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1616 (
  .O(mux_o_1616),
  .I0(ram16s_inst_24_dout[2]),
  .I1(ram16s_inst_25_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1617 (
  .O(mux_o_1617),
  .I0(ram16s_inst_26_dout[2]),
  .I1(ram16s_inst_27_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1618 (
  .O(mux_o_1618),
  .I0(ram16s_inst_28_dout[2]),
  .I1(ram16s_inst_29_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1619 (
  .O(mux_o_1619),
  .I0(ram16s_inst_30_dout[2]),
  .I1(ram16s_inst_31_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1620 (
  .O(mux_o_1620),
  .I0(ram16s_inst_32_dout[2]),
  .I1(ram16s_inst_33_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1621 (
  .O(mux_o_1621),
  .I0(ram16s_inst_34_dout[2]),
  .I1(ram16s_inst_35_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1622 (
  .O(mux_o_1622),
  .I0(ram16s_inst_36_dout[2]),
  .I1(ram16s_inst_37_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1623 (
  .O(mux_o_1623),
  .I0(ram16s_inst_38_dout[2]),
  .I1(ram16s_inst_39_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1624 (
  .O(mux_o_1624),
  .I0(ram16s_inst_40_dout[2]),
  .I1(ram16s_inst_41_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1625 (
  .O(mux_o_1625),
  .I0(ram16s_inst_42_dout[2]),
  .I1(ram16s_inst_43_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1626 (
  .O(mux_o_1626),
  .I0(ram16s_inst_44_dout[2]),
  .I1(ram16s_inst_45_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1627 (
  .O(mux_o_1627),
  .I0(ram16s_inst_46_dout[2]),
  .I1(ram16s_inst_47_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1628 (
  .O(mux_o_1628),
  .I0(ram16s_inst_48_dout[2]),
  .I1(ram16s_inst_49_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1629 (
  .O(mux_o_1629),
  .I0(ram16s_inst_50_dout[2]),
  .I1(ram16s_inst_51_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1630 (
  .O(mux_o_1630),
  .I0(ram16s_inst_52_dout[2]),
  .I1(ram16s_inst_53_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1631 (
  .O(mux_o_1631),
  .I0(ram16s_inst_54_dout[2]),
  .I1(ram16s_inst_55_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1632 (
  .O(mux_o_1632),
  .I0(ram16s_inst_56_dout[2]),
  .I1(ram16s_inst_57_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1633 (
  .O(mux_o_1633),
  .I0(ram16s_inst_58_dout[2]),
  .I1(ram16s_inst_59_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1634 (
  .O(mux_o_1634),
  .I0(ram16s_inst_60_dout[2]),
  .I1(ram16s_inst_61_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1635 (
  .O(mux_o_1635),
  .I0(ram16s_inst_62_dout[2]),
  .I1(ram16s_inst_63_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1636 (
  .O(mux_o_1636),
  .I0(ram16s_inst_64_dout[2]),
  .I1(ram16s_inst_65_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1637 (
  .O(mux_o_1637),
  .I0(ram16s_inst_66_dout[2]),
  .I1(ram16s_inst_67_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1638 (
  .O(mux_o_1638),
  .I0(ram16s_inst_68_dout[2]),
  .I1(ram16s_inst_69_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1639 (
  .O(mux_o_1639),
  .I0(ram16s_inst_70_dout[2]),
  .I1(ram16s_inst_71_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1640 (
  .O(mux_o_1640),
  .I0(ram16s_inst_72_dout[2]),
  .I1(ram16s_inst_73_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1641 (
  .O(mux_o_1641),
  .I0(ram16s_inst_74_dout[2]),
  .I1(ram16s_inst_75_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1642 (
  .O(mux_o_1642),
  .I0(ram16s_inst_76_dout[2]),
  .I1(ram16s_inst_77_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1643 (
  .O(mux_o_1643),
  .I0(ram16s_inst_78_dout[2]),
  .I1(ram16s_inst_79_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1644 (
  .O(mux_o_1644),
  .I0(ram16s_inst_80_dout[2]),
  .I1(ram16s_inst_81_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1645 (
  .O(mux_o_1645),
  .I0(ram16s_inst_82_dout[2]),
  .I1(ram16s_inst_83_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1646 (
  .O(mux_o_1646),
  .I0(ram16s_inst_84_dout[2]),
  .I1(ram16s_inst_85_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1647 (
  .O(mux_o_1647),
  .I0(ram16s_inst_86_dout[2]),
  .I1(ram16s_inst_87_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1648 (
  .O(mux_o_1648),
  .I0(ram16s_inst_88_dout[2]),
  .I1(ram16s_inst_89_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1649 (
  .O(mux_o_1649),
  .I0(ram16s_inst_90_dout[2]),
  .I1(ram16s_inst_91_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1650 (
  .O(mux_o_1650),
  .I0(ram16s_inst_92_dout[2]),
  .I1(ram16s_inst_93_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1651 (
  .O(mux_o_1651),
  .I0(ram16s_inst_94_dout[2]),
  .I1(ram16s_inst_95_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1652 (
  .O(mux_o_1652),
  .I0(ram16s_inst_96_dout[2]),
  .I1(ram16s_inst_97_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1653 (
  .O(mux_o_1653),
  .I0(ram16s_inst_98_dout[2]),
  .I1(ram16s_inst_99_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1654 (
  .O(mux_o_1654),
  .I0(ram16s_inst_100_dout[2]),
  .I1(ram16s_inst_101_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1655 (
  .O(mux_o_1655),
  .I0(ram16s_inst_102_dout[2]),
  .I1(ram16s_inst_103_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1656 (
  .O(mux_o_1656),
  .I0(ram16s_inst_104_dout[2]),
  .I1(ram16s_inst_105_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1657 (
  .O(mux_o_1657),
  .I0(ram16s_inst_106_dout[2]),
  .I1(ram16s_inst_107_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1658 (
  .O(mux_o_1658),
  .I0(ram16s_inst_108_dout[2]),
  .I1(ram16s_inst_109_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1659 (
  .O(mux_o_1659),
  .I0(ram16s_inst_110_dout[2]),
  .I1(ram16s_inst_111_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1660 (
  .O(mux_o_1660),
  .I0(ram16s_inst_112_dout[2]),
  .I1(ram16s_inst_113_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1661 (
  .O(mux_o_1661),
  .I0(ram16s_inst_114_dout[2]),
  .I1(ram16s_inst_115_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1662 (
  .O(mux_o_1662),
  .I0(ram16s_inst_116_dout[2]),
  .I1(ram16s_inst_117_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1663 (
  .O(mux_o_1663),
  .I0(ram16s_inst_118_dout[2]),
  .I1(ram16s_inst_119_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1664 (
  .O(mux_o_1664),
  .I0(ram16s_inst_120_dout[2]),
  .I1(ram16s_inst_121_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1665 (
  .O(mux_o_1665),
  .I0(ram16s_inst_122_dout[2]),
  .I1(ram16s_inst_123_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1666 (
  .O(mux_o_1666),
  .I0(ram16s_inst_124_dout[2]),
  .I1(ram16s_inst_125_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1667 (
  .O(mux_o_1667),
  .I0(ram16s_inst_126_dout[2]),
  .I1(ram16s_inst_127_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1668 (
  .O(mux_o_1668),
  .I0(ram16s_inst_128_dout[2]),
  .I1(ram16s_inst_129_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1669 (
  .O(mux_o_1669),
  .I0(ram16s_inst_130_dout[2]),
  .I1(ram16s_inst_131_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1670 (
  .O(mux_o_1670),
  .I0(ram16s_inst_132_dout[2]),
  .I1(ram16s_inst_133_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1671 (
  .O(mux_o_1671),
  .I0(ram16s_inst_134_dout[2]),
  .I1(ram16s_inst_135_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1672 (
  .O(mux_o_1672),
  .I0(ram16s_inst_136_dout[2]),
  .I1(ram16s_inst_137_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1673 (
  .O(mux_o_1673),
  .I0(ram16s_inst_138_dout[2]),
  .I1(ram16s_inst_139_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1674 (
  .O(mux_o_1674),
  .I0(ram16s_inst_140_dout[2]),
  .I1(ram16s_inst_141_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1675 (
  .O(mux_o_1675),
  .I0(ram16s_inst_142_dout[2]),
  .I1(ram16s_inst_143_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1676 (
  .O(mux_o_1676),
  .I0(ram16s_inst_144_dout[2]),
  .I1(ram16s_inst_145_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1677 (
  .O(mux_o_1677),
  .I0(ram16s_inst_146_dout[2]),
  .I1(ram16s_inst_147_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1678 (
  .O(mux_o_1678),
  .I0(ram16s_inst_148_dout[2]),
  .I1(ram16s_inst_149_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1679 (
  .O(mux_o_1679),
  .I0(ram16s_inst_150_dout[2]),
  .I1(ram16s_inst_151_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1680 (
  .O(mux_o_1680),
  .I0(ram16s_inst_152_dout[2]),
  .I1(ram16s_inst_153_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1681 (
  .O(mux_o_1681),
  .I0(ram16s_inst_154_dout[2]),
  .I1(ram16s_inst_155_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1682 (
  .O(mux_o_1682),
  .I0(ram16s_inst_156_dout[2]),
  .I1(ram16s_inst_157_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1683 (
  .O(mux_o_1683),
  .I0(ram16s_inst_158_dout[2]),
  .I1(ram16s_inst_159_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1684 (
  .O(mux_o_1684),
  .I0(ram16s_inst_160_dout[2]),
  .I1(ram16s_inst_161_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1685 (
  .O(mux_o_1685),
  .I0(ram16s_inst_162_dout[2]),
  .I1(ram16s_inst_163_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1686 (
  .O(mux_o_1686),
  .I0(ram16s_inst_164_dout[2]),
  .I1(ram16s_inst_165_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1687 (
  .O(mux_o_1687),
  .I0(ram16s_inst_166_dout[2]),
  .I1(ram16s_inst_167_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1688 (
  .O(mux_o_1688),
  .I0(ram16s_inst_168_dout[2]),
  .I1(ram16s_inst_169_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1689 (
  .O(mux_o_1689),
  .I0(ram16s_inst_170_dout[2]),
  .I1(ram16s_inst_171_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1690 (
  .O(mux_o_1690),
  .I0(ram16s_inst_172_dout[2]),
  .I1(ram16s_inst_173_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1691 (
  .O(mux_o_1691),
  .I0(ram16s_inst_174_dout[2]),
  .I1(ram16s_inst_175_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1692 (
  .O(mux_o_1692),
  .I0(ram16s_inst_176_dout[2]),
  .I1(ram16s_inst_177_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1693 (
  .O(mux_o_1693),
  .I0(ram16s_inst_178_dout[2]),
  .I1(ram16s_inst_179_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1694 (
  .O(mux_o_1694),
  .I0(ram16s_inst_180_dout[2]),
  .I1(ram16s_inst_181_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1695 (
  .O(mux_o_1695),
  .I0(ram16s_inst_182_dout[2]),
  .I1(ram16s_inst_183_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1696 (
  .O(mux_o_1696),
  .I0(ram16s_inst_184_dout[2]),
  .I1(ram16s_inst_185_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1697 (
  .O(mux_o_1697),
  .I0(ram16s_inst_186_dout[2]),
  .I1(ram16s_inst_187_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1698 (
  .O(mux_o_1698),
  .I0(ram16s_inst_188_dout[2]),
  .I1(ram16s_inst_189_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1699 (
  .O(mux_o_1699),
  .I0(ram16s_inst_190_dout[2]),
  .I1(ram16s_inst_191_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1700 (
  .O(mux_o_1700),
  .I0(ram16s_inst_192_dout[2]),
  .I1(ram16s_inst_193_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1701 (
  .O(mux_o_1701),
  .I0(ram16s_inst_194_dout[2]),
  .I1(ram16s_inst_195_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1702 (
  .O(mux_o_1702),
  .I0(ram16s_inst_196_dout[2]),
  .I1(ram16s_inst_197_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1703 (
  .O(mux_o_1703),
  .I0(ram16s_inst_198_dout[2]),
  .I1(ram16s_inst_199_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1704 (
  .O(mux_o_1704),
  .I0(ram16s_inst_200_dout[2]),
  .I1(ram16s_inst_201_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1705 (
  .O(mux_o_1705),
  .I0(ram16s_inst_202_dout[2]),
  .I1(ram16s_inst_203_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1706 (
  .O(mux_o_1706),
  .I0(ram16s_inst_204_dout[2]),
  .I1(ram16s_inst_205_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1707 (
  .O(mux_o_1707),
  .I0(ram16s_inst_206_dout[2]),
  .I1(ram16s_inst_207_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1708 (
  .O(mux_o_1708),
  .I0(ram16s_inst_208_dout[2]),
  .I1(ram16s_inst_209_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1709 (
  .O(mux_o_1709),
  .I0(ram16s_inst_210_dout[2]),
  .I1(ram16s_inst_211_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1710 (
  .O(mux_o_1710),
  .I0(ram16s_inst_212_dout[2]),
  .I1(ram16s_inst_213_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1711 (
  .O(mux_o_1711),
  .I0(ram16s_inst_214_dout[2]),
  .I1(ram16s_inst_215_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1712 (
  .O(mux_o_1712),
  .I0(ram16s_inst_216_dout[2]),
  .I1(ram16s_inst_217_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1713 (
  .O(mux_o_1713),
  .I0(ram16s_inst_218_dout[2]),
  .I1(ram16s_inst_219_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1714 (
  .O(mux_o_1714),
  .I0(ram16s_inst_220_dout[2]),
  .I1(ram16s_inst_221_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1715 (
  .O(mux_o_1715),
  .I0(ram16s_inst_222_dout[2]),
  .I1(ram16s_inst_223_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1716 (
  .O(mux_o_1716),
  .I0(ram16s_inst_224_dout[2]),
  .I1(ram16s_inst_225_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1717 (
  .O(mux_o_1717),
  .I0(ram16s_inst_226_dout[2]),
  .I1(ram16s_inst_227_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1718 (
  .O(mux_o_1718),
  .I0(ram16s_inst_228_dout[2]),
  .I1(ram16s_inst_229_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1719 (
  .O(mux_o_1719),
  .I0(ram16s_inst_230_dout[2]),
  .I1(ram16s_inst_231_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1720 (
  .O(mux_o_1720),
  .I0(ram16s_inst_232_dout[2]),
  .I1(ram16s_inst_233_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1721 (
  .O(mux_o_1721),
  .I0(ram16s_inst_234_dout[2]),
  .I1(ram16s_inst_235_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1722 (
  .O(mux_o_1722),
  .I0(ram16s_inst_236_dout[2]),
  .I1(ram16s_inst_237_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1723 (
  .O(mux_o_1723),
  .I0(ram16s_inst_238_dout[2]),
  .I1(ram16s_inst_239_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1724 (
  .O(mux_o_1724),
  .I0(ram16s_inst_240_dout[2]),
  .I1(ram16s_inst_241_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1725 (
  .O(mux_o_1725),
  .I0(ram16s_inst_242_dout[2]),
  .I1(ram16s_inst_243_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1726 (
  .O(mux_o_1726),
  .I0(ram16s_inst_244_dout[2]),
  .I1(ram16s_inst_245_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1727 (
  .O(mux_o_1727),
  .I0(ram16s_inst_246_dout[2]),
  .I1(ram16s_inst_247_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1728 (
  .O(mux_o_1728),
  .I0(ram16s_inst_248_dout[2]),
  .I1(ram16s_inst_249_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1729 (
  .O(mux_o_1729),
  .I0(ram16s_inst_250_dout[2]),
  .I1(ram16s_inst_251_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1730 (
  .O(mux_o_1730),
  .I0(ram16s_inst_252_dout[2]),
  .I1(ram16s_inst_253_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1731 (
  .O(mux_o_1731),
  .I0(ram16s_inst_254_dout[2]),
  .I1(ram16s_inst_255_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1732 (
  .O(mux_o_1732),
  .I0(ram16s_inst_256_dout[2]),
  .I1(ram16s_inst_257_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1733 (
  .O(mux_o_1733),
  .I0(ram16s_inst_258_dout[2]),
  .I1(ram16s_inst_259_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1734 (
  .O(mux_o_1734),
  .I0(ram16s_inst_260_dout[2]),
  .I1(ram16s_inst_261_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1735 (
  .O(mux_o_1735),
  .I0(ram16s_inst_262_dout[2]),
  .I1(ram16s_inst_263_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1736 (
  .O(mux_o_1736),
  .I0(ram16s_inst_264_dout[2]),
  .I1(ram16s_inst_265_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1737 (
  .O(mux_o_1737),
  .I0(ram16s_inst_266_dout[2]),
  .I1(ram16s_inst_267_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1738 (
  .O(mux_o_1738),
  .I0(ram16s_inst_268_dout[2]),
  .I1(ram16s_inst_269_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1739 (
  .O(mux_o_1739),
  .I0(ram16s_inst_270_dout[2]),
  .I1(ram16s_inst_271_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1740 (
  .O(mux_o_1740),
  .I0(ram16s_inst_272_dout[2]),
  .I1(ram16s_inst_273_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1741 (
  .O(mux_o_1741),
  .I0(ram16s_inst_274_dout[2]),
  .I1(ram16s_inst_275_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1742 (
  .O(mux_o_1742),
  .I0(ram16s_inst_276_dout[2]),
  .I1(ram16s_inst_277_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1743 (
  .O(mux_o_1743),
  .I0(ram16s_inst_278_dout[2]),
  .I1(ram16s_inst_279_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1744 (
  .O(mux_o_1744),
  .I0(ram16s_inst_280_dout[2]),
  .I1(ram16s_inst_281_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1745 (
  .O(mux_o_1745),
  .I0(ram16s_inst_282_dout[2]),
  .I1(ram16s_inst_283_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1746 (
  .O(mux_o_1746),
  .I0(ram16s_inst_284_dout[2]),
  .I1(ram16s_inst_285_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1747 (
  .O(mux_o_1747),
  .I0(ram16s_inst_286_dout[2]),
  .I1(ram16s_inst_287_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1748 (
  .O(mux_o_1748),
  .I0(ram16s_inst_288_dout[2]),
  .I1(ram16s_inst_289_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1749 (
  .O(mux_o_1749),
  .I0(ram16s_inst_290_dout[2]),
  .I1(ram16s_inst_291_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1750 (
  .O(mux_o_1750),
  .I0(ram16s_inst_292_dout[2]),
  .I1(ram16s_inst_293_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1751 (
  .O(mux_o_1751),
  .I0(ram16s_inst_294_dout[2]),
  .I1(ram16s_inst_295_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1752 (
  .O(mux_o_1752),
  .I0(ram16s_inst_296_dout[2]),
  .I1(ram16s_inst_297_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1753 (
  .O(mux_o_1753),
  .I0(ram16s_inst_298_dout[2]),
  .I1(ram16s_inst_299_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1754 (
  .O(mux_o_1754),
  .I0(ram16s_inst_300_dout[2]),
  .I1(ram16s_inst_301_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1755 (
  .O(mux_o_1755),
  .I0(ram16s_inst_302_dout[2]),
  .I1(ram16s_inst_303_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1756 (
  .O(mux_o_1756),
  .I0(ram16s_inst_304_dout[2]),
  .I1(ram16s_inst_305_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1757 (
  .O(mux_o_1757),
  .I0(ram16s_inst_306_dout[2]),
  .I1(ram16s_inst_307_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1758 (
  .O(mux_o_1758),
  .I0(ram16s_inst_308_dout[2]),
  .I1(ram16s_inst_309_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1759 (
  .O(mux_o_1759),
  .I0(ram16s_inst_310_dout[2]),
  .I1(ram16s_inst_311_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1760 (
  .O(mux_o_1760),
  .I0(ram16s_inst_312_dout[2]),
  .I1(ram16s_inst_313_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1761 (
  .O(mux_o_1761),
  .I0(ram16s_inst_314_dout[2]),
  .I1(ram16s_inst_315_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1762 (
  .O(mux_o_1762),
  .I0(ram16s_inst_316_dout[2]),
  .I1(ram16s_inst_317_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1763 (
  .O(mux_o_1763),
  .I0(ram16s_inst_318_dout[2]),
  .I1(ram16s_inst_319_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1764 (
  .O(mux_o_1764),
  .I0(ram16s_inst_320_dout[2]),
  .I1(ram16s_inst_321_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1765 (
  .O(mux_o_1765),
  .I0(ram16s_inst_322_dout[2]),
  .I1(ram16s_inst_323_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1766 (
  .O(mux_o_1766),
  .I0(ram16s_inst_324_dout[2]),
  .I1(ram16s_inst_325_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1767 (
  .O(mux_o_1767),
  .I0(ram16s_inst_326_dout[2]),
  .I1(ram16s_inst_327_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1768 (
  .O(mux_o_1768),
  .I0(ram16s_inst_328_dout[2]),
  .I1(ram16s_inst_329_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1769 (
  .O(mux_o_1769),
  .I0(ram16s_inst_330_dout[2]),
  .I1(ram16s_inst_331_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1770 (
  .O(mux_o_1770),
  .I0(ram16s_inst_332_dout[2]),
  .I1(ram16s_inst_333_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1771 (
  .O(mux_o_1771),
  .I0(ram16s_inst_334_dout[2]),
  .I1(ram16s_inst_335_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1772 (
  .O(mux_o_1772),
  .I0(ram16s_inst_336_dout[2]),
  .I1(ram16s_inst_337_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1773 (
  .O(mux_o_1773),
  .I0(ram16s_inst_338_dout[2]),
  .I1(ram16s_inst_339_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1774 (
  .O(mux_o_1774),
  .I0(ram16s_inst_340_dout[2]),
  .I1(ram16s_inst_341_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1775 (
  .O(mux_o_1775),
  .I0(ram16s_inst_342_dout[2]),
  .I1(ram16s_inst_343_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1776 (
  .O(mux_o_1776),
  .I0(ram16s_inst_344_dout[2]),
  .I1(ram16s_inst_345_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1777 (
  .O(mux_o_1777),
  .I0(ram16s_inst_346_dout[2]),
  .I1(ram16s_inst_347_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1778 (
  .O(mux_o_1778),
  .I0(ram16s_inst_348_dout[2]),
  .I1(ram16s_inst_349_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1779 (
  .O(mux_o_1779),
  .I0(ram16s_inst_350_dout[2]),
  .I1(ram16s_inst_351_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1780 (
  .O(mux_o_1780),
  .I0(ram16s_inst_352_dout[2]),
  .I1(ram16s_inst_353_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1781 (
  .O(mux_o_1781),
  .I0(ram16s_inst_354_dout[2]),
  .I1(ram16s_inst_355_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1782 (
  .O(mux_o_1782),
  .I0(ram16s_inst_356_dout[2]),
  .I1(ram16s_inst_357_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1783 (
  .O(mux_o_1783),
  .I0(ram16s_inst_358_dout[2]),
  .I1(ram16s_inst_359_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1784 (
  .O(mux_o_1784),
  .I0(ram16s_inst_360_dout[2]),
  .I1(ram16s_inst_361_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1785 (
  .O(mux_o_1785),
  .I0(ram16s_inst_362_dout[2]),
  .I1(ram16s_inst_363_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1786 (
  .O(mux_o_1786),
  .I0(ram16s_inst_364_dout[2]),
  .I1(ram16s_inst_365_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1787 (
  .O(mux_o_1787),
  .I0(ram16s_inst_366_dout[2]),
  .I1(ram16s_inst_367_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1788 (
  .O(mux_o_1788),
  .I0(ram16s_inst_368_dout[2]),
  .I1(ram16s_inst_369_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1789 (
  .O(mux_o_1789),
  .I0(ram16s_inst_370_dout[2]),
  .I1(ram16s_inst_371_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1790 (
  .O(mux_o_1790),
  .I0(ram16s_inst_372_dout[2]),
  .I1(ram16s_inst_373_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1791 (
  .O(mux_o_1791),
  .I0(ram16s_inst_374_dout[2]),
  .I1(ram16s_inst_375_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1792 (
  .O(mux_o_1792),
  .I0(ram16s_inst_376_dout[2]),
  .I1(ram16s_inst_377_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1793 (
  .O(mux_o_1793),
  .I0(ram16s_inst_378_dout[2]),
  .I1(ram16s_inst_379_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1794 (
  .O(mux_o_1794),
  .I0(ram16s_inst_380_dout[2]),
  .I1(ram16s_inst_381_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1795 (
  .O(mux_o_1795),
  .I0(ram16s_inst_382_dout[2]),
  .I1(ram16s_inst_383_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1796 (
  .O(mux_o_1796),
  .I0(ram16s_inst_384_dout[2]),
  .I1(ram16s_inst_385_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1797 (
  .O(mux_o_1797),
  .I0(ram16s_inst_386_dout[2]),
  .I1(ram16s_inst_387_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1798 (
  .O(mux_o_1798),
  .I0(ram16s_inst_388_dout[2]),
  .I1(ram16s_inst_389_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1799 (
  .O(mux_o_1799),
  .I0(ram16s_inst_390_dout[2]),
  .I1(ram16s_inst_391_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1800 (
  .O(mux_o_1800),
  .I0(ram16s_inst_392_dout[2]),
  .I1(ram16s_inst_393_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1801 (
  .O(mux_o_1801),
  .I0(ram16s_inst_394_dout[2]),
  .I1(ram16s_inst_395_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1802 (
  .O(mux_o_1802),
  .I0(ram16s_inst_396_dout[2]),
  .I1(ram16s_inst_397_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1803 (
  .O(mux_o_1803),
  .I0(ram16s_inst_398_dout[2]),
  .I1(ram16s_inst_399_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1804 (
  .O(mux_o_1804),
  .I0(ram16s_inst_400_dout[2]),
  .I1(ram16s_inst_401_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1805 (
  .O(mux_o_1805),
  .I0(ram16s_inst_402_dout[2]),
  .I1(ram16s_inst_403_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1806 (
  .O(mux_o_1806),
  .I0(ram16s_inst_404_dout[2]),
  .I1(ram16s_inst_405_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1807 (
  .O(mux_o_1807),
  .I0(ram16s_inst_406_dout[2]),
  .I1(ram16s_inst_407_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1808 (
  .O(mux_o_1808),
  .I0(ram16s_inst_408_dout[2]),
  .I1(ram16s_inst_409_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1809 (
  .O(mux_o_1809),
  .I0(ram16s_inst_410_dout[2]),
  .I1(ram16s_inst_411_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1810 (
  .O(mux_o_1810),
  .I0(ram16s_inst_412_dout[2]),
  .I1(ram16s_inst_413_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1811 (
  .O(mux_o_1811),
  .I0(ram16s_inst_414_dout[2]),
  .I1(ram16s_inst_415_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1812 (
  .O(mux_o_1812),
  .I0(ram16s_inst_416_dout[2]),
  .I1(ram16s_inst_417_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1813 (
  .O(mux_o_1813),
  .I0(ram16s_inst_418_dout[2]),
  .I1(ram16s_inst_419_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1814 (
  .O(mux_o_1814),
  .I0(ram16s_inst_420_dout[2]),
  .I1(ram16s_inst_421_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1815 (
  .O(mux_o_1815),
  .I0(ram16s_inst_422_dout[2]),
  .I1(ram16s_inst_423_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1816 (
  .O(mux_o_1816),
  .I0(ram16s_inst_424_dout[2]),
  .I1(ram16s_inst_425_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1817 (
  .O(mux_o_1817),
  .I0(ram16s_inst_426_dout[2]),
  .I1(ram16s_inst_427_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1818 (
  .O(mux_o_1818),
  .I0(ram16s_inst_428_dout[2]),
  .I1(ram16s_inst_429_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1819 (
  .O(mux_o_1819),
  .I0(ram16s_inst_430_dout[2]),
  .I1(ram16s_inst_431_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1820 (
  .O(mux_o_1820),
  .I0(ram16s_inst_432_dout[2]),
  .I1(ram16s_inst_433_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1821 (
  .O(mux_o_1821),
  .I0(ram16s_inst_434_dout[2]),
  .I1(ram16s_inst_435_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1822 (
  .O(mux_o_1822),
  .I0(ram16s_inst_436_dout[2]),
  .I1(ram16s_inst_437_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1823 (
  .O(mux_o_1823),
  .I0(ram16s_inst_438_dout[2]),
  .I1(ram16s_inst_439_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1824 (
  .O(mux_o_1824),
  .I0(ram16s_inst_440_dout[2]),
  .I1(ram16s_inst_441_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1825 (
  .O(mux_o_1825),
  .I0(ram16s_inst_442_dout[2]),
  .I1(ram16s_inst_443_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1826 (
  .O(mux_o_1826),
  .I0(ram16s_inst_444_dout[2]),
  .I1(ram16s_inst_445_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1827 (
  .O(mux_o_1827),
  .I0(ram16s_inst_446_dout[2]),
  .I1(ram16s_inst_447_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1828 (
  .O(mux_o_1828),
  .I0(ram16s_inst_448_dout[2]),
  .I1(ram16s_inst_449_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1829 (
  .O(mux_o_1829),
  .I0(ram16s_inst_450_dout[2]),
  .I1(ram16s_inst_451_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1830 (
  .O(mux_o_1830),
  .I0(ram16s_inst_452_dout[2]),
  .I1(ram16s_inst_453_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1831 (
  .O(mux_o_1831),
  .I0(ram16s_inst_454_dout[2]),
  .I1(ram16s_inst_455_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1832 (
  .O(mux_o_1832),
  .I0(ram16s_inst_456_dout[2]),
  .I1(ram16s_inst_457_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1833 (
  .O(mux_o_1833),
  .I0(ram16s_inst_458_dout[2]),
  .I1(ram16s_inst_459_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1834 (
  .O(mux_o_1834),
  .I0(ram16s_inst_460_dout[2]),
  .I1(ram16s_inst_461_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1835 (
  .O(mux_o_1835),
  .I0(ram16s_inst_462_dout[2]),
  .I1(ram16s_inst_463_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1836 (
  .O(mux_o_1836),
  .I0(ram16s_inst_464_dout[2]),
  .I1(ram16s_inst_465_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1837 (
  .O(mux_o_1837),
  .I0(ram16s_inst_466_dout[2]),
  .I1(ram16s_inst_467_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1838 (
  .O(mux_o_1838),
  .I0(ram16s_inst_468_dout[2]),
  .I1(ram16s_inst_469_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1839 (
  .O(mux_o_1839),
  .I0(ram16s_inst_470_dout[2]),
  .I1(ram16s_inst_471_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1840 (
  .O(mux_o_1840),
  .I0(ram16s_inst_472_dout[2]),
  .I1(ram16s_inst_473_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1841 (
  .O(mux_o_1841),
  .I0(ram16s_inst_474_dout[2]),
  .I1(ram16s_inst_475_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1842 (
  .O(mux_o_1842),
  .I0(ram16s_inst_476_dout[2]),
  .I1(ram16s_inst_477_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1843 (
  .O(mux_o_1843),
  .I0(ram16s_inst_478_dout[2]),
  .I1(ram16s_inst_479_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1844 (
  .O(mux_o_1844),
  .I0(ram16s_inst_480_dout[2]),
  .I1(ram16s_inst_481_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1845 (
  .O(mux_o_1845),
  .I0(ram16s_inst_482_dout[2]),
  .I1(ram16s_inst_483_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1846 (
  .O(mux_o_1846),
  .I0(ram16s_inst_484_dout[2]),
  .I1(ram16s_inst_485_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1847 (
  .O(mux_o_1847),
  .I0(ram16s_inst_486_dout[2]),
  .I1(ram16s_inst_487_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1848 (
  .O(mux_o_1848),
  .I0(ram16s_inst_488_dout[2]),
  .I1(ram16s_inst_489_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1849 (
  .O(mux_o_1849),
  .I0(ram16s_inst_490_dout[2]),
  .I1(ram16s_inst_491_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1850 (
  .O(mux_o_1850),
  .I0(ram16s_inst_492_dout[2]),
  .I1(ram16s_inst_493_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1851 (
  .O(mux_o_1851),
  .I0(ram16s_inst_494_dout[2]),
  .I1(ram16s_inst_495_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1852 (
  .O(mux_o_1852),
  .I0(ram16s_inst_496_dout[2]),
  .I1(ram16s_inst_497_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1853 (
  .O(mux_o_1853),
  .I0(ram16s_inst_498_dout[2]),
  .I1(ram16s_inst_499_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1854 (
  .O(mux_o_1854),
  .I0(ram16s_inst_500_dout[2]),
  .I1(ram16s_inst_501_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1855 (
  .O(mux_o_1855),
  .I0(ram16s_inst_502_dout[2]),
  .I1(ram16s_inst_503_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1856 (
  .O(mux_o_1856),
  .I0(ram16s_inst_504_dout[2]),
  .I1(ram16s_inst_505_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1857 (
  .O(mux_o_1857),
  .I0(ram16s_inst_506_dout[2]),
  .I1(ram16s_inst_507_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1858 (
  .O(mux_o_1858),
  .I0(ram16s_inst_508_dout[2]),
  .I1(ram16s_inst_509_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1859 (
  .O(mux_o_1859),
  .I0(ram16s_inst_510_dout[2]),
  .I1(ram16s_inst_511_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1860 (
  .O(mux_o_1860),
  .I0(ram16s_inst_512_dout[2]),
  .I1(ram16s_inst_513_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1861 (
  .O(mux_o_1861),
  .I0(ram16s_inst_514_dout[2]),
  .I1(ram16s_inst_515_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1862 (
  .O(mux_o_1862),
  .I0(ram16s_inst_516_dout[2]),
  .I1(ram16s_inst_517_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1863 (
  .O(mux_o_1863),
  .I0(ram16s_inst_518_dout[2]),
  .I1(ram16s_inst_519_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1864 (
  .O(mux_o_1864),
  .I0(ram16s_inst_520_dout[2]),
  .I1(ram16s_inst_521_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1865 (
  .O(mux_o_1865),
  .I0(ram16s_inst_522_dout[2]),
  .I1(ram16s_inst_523_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1866 (
  .O(mux_o_1866),
  .I0(ram16s_inst_524_dout[2]),
  .I1(ram16s_inst_525_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1867 (
  .O(mux_o_1867),
  .I0(ram16s_inst_526_dout[2]),
  .I1(ram16s_inst_527_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1868 (
  .O(mux_o_1868),
  .I0(ram16s_inst_528_dout[2]),
  .I1(ram16s_inst_529_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1869 (
  .O(mux_o_1869),
  .I0(ram16s_inst_530_dout[2]),
  .I1(ram16s_inst_531_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1870 (
  .O(mux_o_1870),
  .I0(ram16s_inst_532_dout[2]),
  .I1(ram16s_inst_533_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1871 (
  .O(mux_o_1871),
  .I0(ram16s_inst_534_dout[2]),
  .I1(ram16s_inst_535_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1872 (
  .O(mux_o_1872),
  .I0(ram16s_inst_536_dout[2]),
  .I1(ram16s_inst_537_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1873 (
  .O(mux_o_1873),
  .I0(ram16s_inst_538_dout[2]),
  .I1(ram16s_inst_539_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1874 (
  .O(mux_o_1874),
  .I0(ram16s_inst_540_dout[2]),
  .I1(ram16s_inst_541_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1875 (
  .O(mux_o_1875),
  .I0(ram16s_inst_542_dout[2]),
  .I1(ram16s_inst_543_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1876 (
  .O(mux_o_1876),
  .I0(ram16s_inst_544_dout[2]),
  .I1(ram16s_inst_545_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1877 (
  .O(mux_o_1877),
  .I0(ram16s_inst_546_dout[2]),
  .I1(ram16s_inst_547_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1878 (
  .O(mux_o_1878),
  .I0(ram16s_inst_548_dout[2]),
  .I1(ram16s_inst_549_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1879 (
  .O(mux_o_1879),
  .I0(ram16s_inst_550_dout[2]),
  .I1(ram16s_inst_551_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1880 (
  .O(mux_o_1880),
  .I0(ram16s_inst_552_dout[2]),
  .I1(ram16s_inst_553_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1881 (
  .O(mux_o_1881),
  .I0(ram16s_inst_554_dout[2]),
  .I1(ram16s_inst_555_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1882 (
  .O(mux_o_1882),
  .I0(ram16s_inst_556_dout[2]),
  .I1(ram16s_inst_557_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1883 (
  .O(mux_o_1883),
  .I0(ram16s_inst_558_dout[2]),
  .I1(ram16s_inst_559_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1884 (
  .O(mux_o_1884),
  .I0(ram16s_inst_560_dout[2]),
  .I1(ram16s_inst_561_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1885 (
  .O(mux_o_1885),
  .I0(ram16s_inst_562_dout[2]),
  .I1(ram16s_inst_563_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1886 (
  .O(mux_o_1886),
  .I0(ram16s_inst_564_dout[2]),
  .I1(ram16s_inst_565_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1887 (
  .O(mux_o_1887),
  .I0(ram16s_inst_566_dout[2]),
  .I1(ram16s_inst_567_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1888 (
  .O(mux_o_1888),
  .I0(ram16s_inst_568_dout[2]),
  .I1(ram16s_inst_569_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1889 (
  .O(mux_o_1889),
  .I0(ram16s_inst_570_dout[2]),
  .I1(ram16s_inst_571_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1890 (
  .O(mux_o_1890),
  .I0(ram16s_inst_572_dout[2]),
  .I1(ram16s_inst_573_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1891 (
  .O(mux_o_1891),
  .I0(ram16s_inst_574_dout[2]),
  .I1(ram16s_inst_575_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1892 (
  .O(mux_o_1892),
  .I0(ram16s_inst_576_dout[2]),
  .I1(ram16s_inst_577_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1893 (
  .O(mux_o_1893),
  .I0(ram16s_inst_578_dout[2]),
  .I1(ram16s_inst_579_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1894 (
  .O(mux_o_1894),
  .I0(ram16s_inst_580_dout[2]),
  .I1(ram16s_inst_581_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1895 (
  .O(mux_o_1895),
  .I0(ram16s_inst_582_dout[2]),
  .I1(ram16s_inst_583_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1896 (
  .O(mux_o_1896),
  .I0(ram16s_inst_584_dout[2]),
  .I1(ram16s_inst_585_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1897 (
  .O(mux_o_1897),
  .I0(ram16s_inst_586_dout[2]),
  .I1(ram16s_inst_587_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1898 (
  .O(mux_o_1898),
  .I0(ram16s_inst_588_dout[2]),
  .I1(ram16s_inst_589_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1899 (
  .O(mux_o_1899),
  .I0(ram16s_inst_590_dout[2]),
  .I1(ram16s_inst_591_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1900 (
  .O(mux_o_1900),
  .I0(ram16s_inst_592_dout[2]),
  .I1(ram16s_inst_593_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1901 (
  .O(mux_o_1901),
  .I0(ram16s_inst_594_dout[2]),
  .I1(ram16s_inst_595_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1902 (
  .O(mux_o_1902),
  .I0(ram16s_inst_596_dout[2]),
  .I1(ram16s_inst_597_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1903 (
  .O(mux_o_1903),
  .I0(ram16s_inst_598_dout[2]),
  .I1(ram16s_inst_599_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1904 (
  .O(mux_o_1904),
  .I0(ram16s_inst_600_dout[2]),
  .I1(ram16s_inst_601_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1905 (
  .O(mux_o_1905),
  .I0(ram16s_inst_602_dout[2]),
  .I1(ram16s_inst_603_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1906 (
  .O(mux_o_1906),
  .I0(ram16s_inst_604_dout[2]),
  .I1(ram16s_inst_605_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1907 (
  .O(mux_o_1907),
  .I0(ram16s_inst_606_dout[2]),
  .I1(ram16s_inst_607_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1908 (
  .O(mux_o_1908),
  .I0(ram16s_inst_608_dout[2]),
  .I1(ram16s_inst_609_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1909 (
  .O(mux_o_1909),
  .I0(ram16s_inst_610_dout[2]),
  .I1(ram16s_inst_611_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1910 (
  .O(mux_o_1910),
  .I0(ram16s_inst_612_dout[2]),
  .I1(ram16s_inst_613_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1911 (
  .O(mux_o_1911),
  .I0(ram16s_inst_614_dout[2]),
  .I1(ram16s_inst_615_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1912 (
  .O(mux_o_1912),
  .I0(ram16s_inst_616_dout[2]),
  .I1(ram16s_inst_617_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1913 (
  .O(mux_o_1913),
  .I0(ram16s_inst_618_dout[2]),
  .I1(ram16s_inst_619_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1914 (
  .O(mux_o_1914),
  .I0(ram16s_inst_620_dout[2]),
  .I1(ram16s_inst_621_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1915 (
  .O(mux_o_1915),
  .I0(ram16s_inst_622_dout[2]),
  .I1(ram16s_inst_623_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1916 (
  .O(mux_o_1916),
  .I0(ram16s_inst_624_dout[2]),
  .I1(ram16s_inst_625_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1917 (
  .O(mux_o_1917),
  .I0(ram16s_inst_626_dout[2]),
  .I1(ram16s_inst_627_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1918 (
  .O(mux_o_1918),
  .I0(ram16s_inst_628_dout[2]),
  .I1(ram16s_inst_629_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1919 (
  .O(mux_o_1919),
  .I0(ram16s_inst_630_dout[2]),
  .I1(ram16s_inst_631_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1920 (
  .O(mux_o_1920),
  .I0(ram16s_inst_632_dout[2]),
  .I1(ram16s_inst_633_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1921 (
  .O(mux_o_1921),
  .I0(ram16s_inst_634_dout[2]),
  .I1(ram16s_inst_635_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1922 (
  .O(mux_o_1922),
  .I0(ram16s_inst_636_dout[2]),
  .I1(ram16s_inst_637_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1923 (
  .O(mux_o_1923),
  .I0(ram16s_inst_638_dout[2]),
  .I1(ram16s_inst_639_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1924 (
  .O(mux_o_1924),
  .I0(ram16s_inst_640_dout[2]),
  .I1(ram16s_inst_641_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1925 (
  .O(mux_o_1925),
  .I0(ram16s_inst_642_dout[2]),
  .I1(ram16s_inst_643_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1926 (
  .O(mux_o_1926),
  .I0(ram16s_inst_644_dout[2]),
  .I1(ram16s_inst_645_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1927 (
  .O(mux_o_1927),
  .I0(ram16s_inst_646_dout[2]),
  .I1(ram16s_inst_647_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1928 (
  .O(mux_o_1928),
  .I0(ram16s_inst_648_dout[2]),
  .I1(ram16s_inst_649_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1929 (
  .O(mux_o_1929),
  .I0(ram16s_inst_650_dout[2]),
  .I1(ram16s_inst_651_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1930 (
  .O(mux_o_1930),
  .I0(ram16s_inst_652_dout[2]),
  .I1(ram16s_inst_653_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1931 (
  .O(mux_o_1931),
  .I0(ram16s_inst_654_dout[2]),
  .I1(ram16s_inst_655_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1932 (
  .O(mux_o_1932),
  .I0(ram16s_inst_656_dout[2]),
  .I1(ram16s_inst_657_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1933 (
  .O(mux_o_1933),
  .I0(ram16s_inst_658_dout[2]),
  .I1(ram16s_inst_659_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1934 (
  .O(mux_o_1934),
  .I0(ram16s_inst_660_dout[2]),
  .I1(ram16s_inst_661_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1935 (
  .O(mux_o_1935),
  .I0(ram16s_inst_662_dout[2]),
  .I1(ram16s_inst_663_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1936 (
  .O(mux_o_1936),
  .I0(ram16s_inst_664_dout[2]),
  .I1(ram16s_inst_665_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1937 (
  .O(mux_o_1937),
  .I0(ram16s_inst_666_dout[2]),
  .I1(ram16s_inst_667_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1938 (
  .O(mux_o_1938),
  .I0(ram16s_inst_668_dout[2]),
  .I1(ram16s_inst_669_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1939 (
  .O(mux_o_1939),
  .I0(ram16s_inst_670_dout[2]),
  .I1(ram16s_inst_671_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1940 (
  .O(mux_o_1940),
  .I0(ram16s_inst_672_dout[2]),
  .I1(ram16s_inst_673_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1941 (
  .O(mux_o_1941),
  .I0(ram16s_inst_674_dout[2]),
  .I1(ram16s_inst_675_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1942 (
  .O(mux_o_1942),
  .I0(ram16s_inst_676_dout[2]),
  .I1(ram16s_inst_677_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1943 (
  .O(mux_o_1943),
  .I0(ram16s_inst_678_dout[2]),
  .I1(ram16s_inst_679_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1944 (
  .O(mux_o_1944),
  .I0(ram16s_inst_680_dout[2]),
  .I1(ram16s_inst_681_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1945 (
  .O(mux_o_1945),
  .I0(ram16s_inst_682_dout[2]),
  .I1(ram16s_inst_683_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1946 (
  .O(mux_o_1946),
  .I0(ram16s_inst_684_dout[2]),
  .I1(ram16s_inst_685_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1947 (
  .O(mux_o_1947),
  .I0(ram16s_inst_686_dout[2]),
  .I1(ram16s_inst_687_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1948 (
  .O(mux_o_1948),
  .I0(ram16s_inst_688_dout[2]),
  .I1(ram16s_inst_689_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1949 (
  .O(mux_o_1949),
  .I0(ram16s_inst_690_dout[2]),
  .I1(ram16s_inst_691_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1950 (
  .O(mux_o_1950),
  .I0(ram16s_inst_692_dout[2]),
  .I1(ram16s_inst_693_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1951 (
  .O(mux_o_1951),
  .I0(ram16s_inst_694_dout[2]),
  .I1(ram16s_inst_695_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1952 (
  .O(mux_o_1952),
  .I0(ram16s_inst_696_dout[2]),
  .I1(ram16s_inst_697_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1953 (
  .O(mux_o_1953),
  .I0(ram16s_inst_698_dout[2]),
  .I1(ram16s_inst_699_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1954 (
  .O(mux_o_1954),
  .I0(ram16s_inst_700_dout[2]),
  .I1(ram16s_inst_701_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1955 (
  .O(mux_o_1955),
  .I0(ram16s_inst_702_dout[2]),
  .I1(ram16s_inst_703_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1956 (
  .O(mux_o_1956),
  .I0(ram16s_inst_704_dout[2]),
  .I1(ram16s_inst_705_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1957 (
  .O(mux_o_1957),
  .I0(ram16s_inst_706_dout[2]),
  .I1(ram16s_inst_707_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1958 (
  .O(mux_o_1958),
  .I0(ram16s_inst_708_dout[2]),
  .I1(ram16s_inst_709_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1959 (
  .O(mux_o_1959),
  .I0(ram16s_inst_710_dout[2]),
  .I1(ram16s_inst_711_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1960 (
  .O(mux_o_1960),
  .I0(ram16s_inst_712_dout[2]),
  .I1(ram16s_inst_713_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1961 (
  .O(mux_o_1961),
  .I0(ram16s_inst_714_dout[2]),
  .I1(ram16s_inst_715_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1962 (
  .O(mux_o_1962),
  .I0(ram16s_inst_716_dout[2]),
  .I1(ram16s_inst_717_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1963 (
  .O(mux_o_1963),
  .I0(ram16s_inst_718_dout[2]),
  .I1(ram16s_inst_719_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1964 (
  .O(mux_o_1964),
  .I0(ram16s_inst_720_dout[2]),
  .I1(ram16s_inst_721_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1965 (
  .O(mux_o_1965),
  .I0(ram16s_inst_722_dout[2]),
  .I1(ram16s_inst_723_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1966 (
  .O(mux_o_1966),
  .I0(ram16s_inst_724_dout[2]),
  .I1(ram16s_inst_725_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1967 (
  .O(mux_o_1967),
  .I0(ram16s_inst_726_dout[2]),
  .I1(ram16s_inst_727_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1968 (
  .O(mux_o_1968),
  .I0(ram16s_inst_728_dout[2]),
  .I1(ram16s_inst_729_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1969 (
  .O(mux_o_1969),
  .I0(ram16s_inst_730_dout[2]),
  .I1(ram16s_inst_731_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1970 (
  .O(mux_o_1970),
  .I0(ram16s_inst_732_dout[2]),
  .I1(ram16s_inst_733_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1971 (
  .O(mux_o_1971),
  .I0(ram16s_inst_734_dout[2]),
  .I1(ram16s_inst_735_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1972 (
  .O(mux_o_1972),
  .I0(ram16s_inst_736_dout[2]),
  .I1(ram16s_inst_737_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1973 (
  .O(mux_o_1973),
  .I0(ram16s_inst_738_dout[2]),
  .I1(ram16s_inst_739_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1974 (
  .O(mux_o_1974),
  .I0(ram16s_inst_740_dout[2]),
  .I1(ram16s_inst_741_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1975 (
  .O(mux_o_1975),
  .I0(ram16s_inst_742_dout[2]),
  .I1(ram16s_inst_743_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1976 (
  .O(mux_o_1976),
  .I0(ram16s_inst_744_dout[2]),
  .I1(ram16s_inst_745_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1977 (
  .O(mux_o_1977),
  .I0(ram16s_inst_746_dout[2]),
  .I1(ram16s_inst_747_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1978 (
  .O(mux_o_1978),
  .I0(ram16s_inst_748_dout[2]),
  .I1(ram16s_inst_749_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1979 (
  .O(mux_o_1979),
  .I0(ram16s_inst_750_dout[2]),
  .I1(ram16s_inst_751_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1980 (
  .O(mux_o_1980),
  .I0(ram16s_inst_752_dout[2]),
  .I1(ram16s_inst_753_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1981 (
  .O(mux_o_1981),
  .I0(ram16s_inst_754_dout[2]),
  .I1(ram16s_inst_755_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1982 (
  .O(mux_o_1982),
  .I0(ram16s_inst_756_dout[2]),
  .I1(ram16s_inst_757_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1983 (
  .O(mux_o_1983),
  .I0(ram16s_inst_758_dout[2]),
  .I1(ram16s_inst_759_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1984 (
  .O(mux_o_1984),
  .I0(ram16s_inst_760_dout[2]),
  .I1(ram16s_inst_761_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1985 (
  .O(mux_o_1985),
  .I0(ram16s_inst_762_dout[2]),
  .I1(ram16s_inst_763_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1986 (
  .O(mux_o_1986),
  .I0(ram16s_inst_764_dout[2]),
  .I1(ram16s_inst_765_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1987 (
  .O(mux_o_1987),
  .I0(ram16s_inst_766_dout[2]),
  .I1(ram16s_inst_767_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1988 (
  .O(mux_o_1988),
  .I0(ram16s_inst_768_dout[2]),
  .I1(ram16s_inst_769_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1989 (
  .O(mux_o_1989),
  .I0(ram16s_inst_770_dout[2]),
  .I1(ram16s_inst_771_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1990 (
  .O(mux_o_1990),
  .I0(ram16s_inst_772_dout[2]),
  .I1(ram16s_inst_773_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1991 (
  .O(mux_o_1991),
  .I0(ram16s_inst_774_dout[2]),
  .I1(ram16s_inst_775_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1992 (
  .O(mux_o_1992),
  .I0(ram16s_inst_776_dout[2]),
  .I1(ram16s_inst_777_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1993 (
  .O(mux_o_1993),
  .I0(ram16s_inst_778_dout[2]),
  .I1(ram16s_inst_779_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1994 (
  .O(mux_o_1994),
  .I0(ram16s_inst_780_dout[2]),
  .I1(ram16s_inst_781_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1995 (
  .O(mux_o_1995),
  .I0(ram16s_inst_782_dout[2]),
  .I1(ram16s_inst_783_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1996 (
  .O(mux_o_1996),
  .I0(ram16s_inst_784_dout[2]),
  .I1(ram16s_inst_785_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1997 (
  .O(mux_o_1997),
  .I0(ram16s_inst_786_dout[2]),
  .I1(ram16s_inst_787_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1998 (
  .O(mux_o_1998),
  .I0(ram16s_inst_788_dout[2]),
  .I1(ram16s_inst_789_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_1999 (
  .O(mux_o_1999),
  .I0(ram16s_inst_790_dout[2]),
  .I1(ram16s_inst_791_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_2000 (
  .O(mux_o_2000),
  .I0(ram16s_inst_792_dout[2]),
  .I1(ram16s_inst_793_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_2001 (
  .O(mux_o_2001),
  .I0(ram16s_inst_794_dout[2]),
  .I1(ram16s_inst_795_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_2002 (
  .O(mux_o_2002),
  .I0(ram16s_inst_796_dout[2]),
  .I1(ram16s_inst_797_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_2003 (
  .O(mux_o_2003),
  .I0(ram16s_inst_798_dout[2]),
  .I1(ram16s_inst_799_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_2004 (
  .O(mux_o_2004),
  .I0(mux_o_1604),
  .I1(mux_o_1605),
  .S0(ad[5])
);
MUX2 mux_inst_2005 (
  .O(mux_o_2005),
  .I0(mux_o_1606),
  .I1(mux_o_1607),
  .S0(ad[5])
);
MUX2 mux_inst_2006 (
  .O(mux_o_2006),
  .I0(mux_o_1608),
  .I1(mux_o_1609),
  .S0(ad[5])
);
MUX2 mux_inst_2007 (
  .O(mux_o_2007),
  .I0(mux_o_1610),
  .I1(mux_o_1611),
  .S0(ad[5])
);
MUX2 mux_inst_2008 (
  .O(mux_o_2008),
  .I0(mux_o_1612),
  .I1(mux_o_1613),
  .S0(ad[5])
);
MUX2 mux_inst_2009 (
  .O(mux_o_2009),
  .I0(mux_o_1614),
  .I1(mux_o_1615),
  .S0(ad[5])
);
MUX2 mux_inst_2010 (
  .O(mux_o_2010),
  .I0(mux_o_1616),
  .I1(mux_o_1617),
  .S0(ad[5])
);
MUX2 mux_inst_2011 (
  .O(mux_o_2011),
  .I0(mux_o_1618),
  .I1(mux_o_1619),
  .S0(ad[5])
);
MUX2 mux_inst_2012 (
  .O(mux_o_2012),
  .I0(mux_o_1620),
  .I1(mux_o_1621),
  .S0(ad[5])
);
MUX2 mux_inst_2013 (
  .O(mux_o_2013),
  .I0(mux_o_1622),
  .I1(mux_o_1623),
  .S0(ad[5])
);
MUX2 mux_inst_2014 (
  .O(mux_o_2014),
  .I0(mux_o_1624),
  .I1(mux_o_1625),
  .S0(ad[5])
);
MUX2 mux_inst_2015 (
  .O(mux_o_2015),
  .I0(mux_o_1626),
  .I1(mux_o_1627),
  .S0(ad[5])
);
MUX2 mux_inst_2016 (
  .O(mux_o_2016),
  .I0(mux_o_1628),
  .I1(mux_o_1629),
  .S0(ad[5])
);
MUX2 mux_inst_2017 (
  .O(mux_o_2017),
  .I0(mux_o_1630),
  .I1(mux_o_1631),
  .S0(ad[5])
);
MUX2 mux_inst_2018 (
  .O(mux_o_2018),
  .I0(mux_o_1632),
  .I1(mux_o_1633),
  .S0(ad[5])
);
MUX2 mux_inst_2019 (
  .O(mux_o_2019),
  .I0(mux_o_1634),
  .I1(mux_o_1635),
  .S0(ad[5])
);
MUX2 mux_inst_2020 (
  .O(mux_o_2020),
  .I0(mux_o_1636),
  .I1(mux_o_1637),
  .S0(ad[5])
);
MUX2 mux_inst_2021 (
  .O(mux_o_2021),
  .I0(mux_o_1638),
  .I1(mux_o_1639),
  .S0(ad[5])
);
MUX2 mux_inst_2022 (
  .O(mux_o_2022),
  .I0(mux_o_1640),
  .I1(mux_o_1641),
  .S0(ad[5])
);
MUX2 mux_inst_2023 (
  .O(mux_o_2023),
  .I0(mux_o_1642),
  .I1(mux_o_1643),
  .S0(ad[5])
);
MUX2 mux_inst_2024 (
  .O(mux_o_2024),
  .I0(mux_o_1644),
  .I1(mux_o_1645),
  .S0(ad[5])
);
MUX2 mux_inst_2025 (
  .O(mux_o_2025),
  .I0(mux_o_1646),
  .I1(mux_o_1647),
  .S0(ad[5])
);
MUX2 mux_inst_2026 (
  .O(mux_o_2026),
  .I0(mux_o_1648),
  .I1(mux_o_1649),
  .S0(ad[5])
);
MUX2 mux_inst_2027 (
  .O(mux_o_2027),
  .I0(mux_o_1650),
  .I1(mux_o_1651),
  .S0(ad[5])
);
MUX2 mux_inst_2028 (
  .O(mux_o_2028),
  .I0(mux_o_1652),
  .I1(mux_o_1653),
  .S0(ad[5])
);
MUX2 mux_inst_2029 (
  .O(mux_o_2029),
  .I0(mux_o_1654),
  .I1(mux_o_1655),
  .S0(ad[5])
);
MUX2 mux_inst_2030 (
  .O(mux_o_2030),
  .I0(mux_o_1656),
  .I1(mux_o_1657),
  .S0(ad[5])
);
MUX2 mux_inst_2031 (
  .O(mux_o_2031),
  .I0(mux_o_1658),
  .I1(mux_o_1659),
  .S0(ad[5])
);
MUX2 mux_inst_2032 (
  .O(mux_o_2032),
  .I0(mux_o_1660),
  .I1(mux_o_1661),
  .S0(ad[5])
);
MUX2 mux_inst_2033 (
  .O(mux_o_2033),
  .I0(mux_o_1662),
  .I1(mux_o_1663),
  .S0(ad[5])
);
MUX2 mux_inst_2034 (
  .O(mux_o_2034),
  .I0(mux_o_1664),
  .I1(mux_o_1665),
  .S0(ad[5])
);
MUX2 mux_inst_2035 (
  .O(mux_o_2035),
  .I0(mux_o_1666),
  .I1(mux_o_1667),
  .S0(ad[5])
);
MUX2 mux_inst_2036 (
  .O(mux_o_2036),
  .I0(mux_o_1668),
  .I1(mux_o_1669),
  .S0(ad[5])
);
MUX2 mux_inst_2037 (
  .O(mux_o_2037),
  .I0(mux_o_1670),
  .I1(mux_o_1671),
  .S0(ad[5])
);
MUX2 mux_inst_2038 (
  .O(mux_o_2038),
  .I0(mux_o_1672),
  .I1(mux_o_1673),
  .S0(ad[5])
);
MUX2 mux_inst_2039 (
  .O(mux_o_2039),
  .I0(mux_o_1674),
  .I1(mux_o_1675),
  .S0(ad[5])
);
MUX2 mux_inst_2040 (
  .O(mux_o_2040),
  .I0(mux_o_1676),
  .I1(mux_o_1677),
  .S0(ad[5])
);
MUX2 mux_inst_2041 (
  .O(mux_o_2041),
  .I0(mux_o_1678),
  .I1(mux_o_1679),
  .S0(ad[5])
);
MUX2 mux_inst_2042 (
  .O(mux_o_2042),
  .I0(mux_o_1680),
  .I1(mux_o_1681),
  .S0(ad[5])
);
MUX2 mux_inst_2043 (
  .O(mux_o_2043),
  .I0(mux_o_1682),
  .I1(mux_o_1683),
  .S0(ad[5])
);
MUX2 mux_inst_2044 (
  .O(mux_o_2044),
  .I0(mux_o_1684),
  .I1(mux_o_1685),
  .S0(ad[5])
);
MUX2 mux_inst_2045 (
  .O(mux_o_2045),
  .I0(mux_o_1686),
  .I1(mux_o_1687),
  .S0(ad[5])
);
MUX2 mux_inst_2046 (
  .O(mux_o_2046),
  .I0(mux_o_1688),
  .I1(mux_o_1689),
  .S0(ad[5])
);
MUX2 mux_inst_2047 (
  .O(mux_o_2047),
  .I0(mux_o_1690),
  .I1(mux_o_1691),
  .S0(ad[5])
);
MUX2 mux_inst_2048 (
  .O(mux_o_2048),
  .I0(mux_o_1692),
  .I1(mux_o_1693),
  .S0(ad[5])
);
MUX2 mux_inst_2049 (
  .O(mux_o_2049),
  .I0(mux_o_1694),
  .I1(mux_o_1695),
  .S0(ad[5])
);
MUX2 mux_inst_2050 (
  .O(mux_o_2050),
  .I0(mux_o_1696),
  .I1(mux_o_1697),
  .S0(ad[5])
);
MUX2 mux_inst_2051 (
  .O(mux_o_2051),
  .I0(mux_o_1698),
  .I1(mux_o_1699),
  .S0(ad[5])
);
MUX2 mux_inst_2052 (
  .O(mux_o_2052),
  .I0(mux_o_1700),
  .I1(mux_o_1701),
  .S0(ad[5])
);
MUX2 mux_inst_2053 (
  .O(mux_o_2053),
  .I0(mux_o_1702),
  .I1(mux_o_1703),
  .S0(ad[5])
);
MUX2 mux_inst_2054 (
  .O(mux_o_2054),
  .I0(mux_o_1704),
  .I1(mux_o_1705),
  .S0(ad[5])
);
MUX2 mux_inst_2055 (
  .O(mux_o_2055),
  .I0(mux_o_1706),
  .I1(mux_o_1707),
  .S0(ad[5])
);
MUX2 mux_inst_2056 (
  .O(mux_o_2056),
  .I0(mux_o_1708),
  .I1(mux_o_1709),
  .S0(ad[5])
);
MUX2 mux_inst_2057 (
  .O(mux_o_2057),
  .I0(mux_o_1710),
  .I1(mux_o_1711),
  .S0(ad[5])
);
MUX2 mux_inst_2058 (
  .O(mux_o_2058),
  .I0(mux_o_1712),
  .I1(mux_o_1713),
  .S0(ad[5])
);
MUX2 mux_inst_2059 (
  .O(mux_o_2059),
  .I0(mux_o_1714),
  .I1(mux_o_1715),
  .S0(ad[5])
);
MUX2 mux_inst_2060 (
  .O(mux_o_2060),
  .I0(mux_o_1716),
  .I1(mux_o_1717),
  .S0(ad[5])
);
MUX2 mux_inst_2061 (
  .O(mux_o_2061),
  .I0(mux_o_1718),
  .I1(mux_o_1719),
  .S0(ad[5])
);
MUX2 mux_inst_2062 (
  .O(mux_o_2062),
  .I0(mux_o_1720),
  .I1(mux_o_1721),
  .S0(ad[5])
);
MUX2 mux_inst_2063 (
  .O(mux_o_2063),
  .I0(mux_o_1722),
  .I1(mux_o_1723),
  .S0(ad[5])
);
MUX2 mux_inst_2064 (
  .O(mux_o_2064),
  .I0(mux_o_1724),
  .I1(mux_o_1725),
  .S0(ad[5])
);
MUX2 mux_inst_2065 (
  .O(mux_o_2065),
  .I0(mux_o_1726),
  .I1(mux_o_1727),
  .S0(ad[5])
);
MUX2 mux_inst_2066 (
  .O(mux_o_2066),
  .I0(mux_o_1728),
  .I1(mux_o_1729),
  .S0(ad[5])
);
MUX2 mux_inst_2067 (
  .O(mux_o_2067),
  .I0(mux_o_1730),
  .I1(mux_o_1731),
  .S0(ad[5])
);
MUX2 mux_inst_2068 (
  .O(mux_o_2068),
  .I0(mux_o_1732),
  .I1(mux_o_1733),
  .S0(ad[5])
);
MUX2 mux_inst_2069 (
  .O(mux_o_2069),
  .I0(mux_o_1734),
  .I1(mux_o_1735),
  .S0(ad[5])
);
MUX2 mux_inst_2070 (
  .O(mux_o_2070),
  .I0(mux_o_1736),
  .I1(mux_o_1737),
  .S0(ad[5])
);
MUX2 mux_inst_2071 (
  .O(mux_o_2071),
  .I0(mux_o_1738),
  .I1(mux_o_1739),
  .S0(ad[5])
);
MUX2 mux_inst_2072 (
  .O(mux_o_2072),
  .I0(mux_o_1740),
  .I1(mux_o_1741),
  .S0(ad[5])
);
MUX2 mux_inst_2073 (
  .O(mux_o_2073),
  .I0(mux_o_1742),
  .I1(mux_o_1743),
  .S0(ad[5])
);
MUX2 mux_inst_2074 (
  .O(mux_o_2074),
  .I0(mux_o_1744),
  .I1(mux_o_1745),
  .S0(ad[5])
);
MUX2 mux_inst_2075 (
  .O(mux_o_2075),
  .I0(mux_o_1746),
  .I1(mux_o_1747),
  .S0(ad[5])
);
MUX2 mux_inst_2076 (
  .O(mux_o_2076),
  .I0(mux_o_1748),
  .I1(mux_o_1749),
  .S0(ad[5])
);
MUX2 mux_inst_2077 (
  .O(mux_o_2077),
  .I0(mux_o_1750),
  .I1(mux_o_1751),
  .S0(ad[5])
);
MUX2 mux_inst_2078 (
  .O(mux_o_2078),
  .I0(mux_o_1752),
  .I1(mux_o_1753),
  .S0(ad[5])
);
MUX2 mux_inst_2079 (
  .O(mux_o_2079),
  .I0(mux_o_1754),
  .I1(mux_o_1755),
  .S0(ad[5])
);
MUX2 mux_inst_2080 (
  .O(mux_o_2080),
  .I0(mux_o_1756),
  .I1(mux_o_1757),
  .S0(ad[5])
);
MUX2 mux_inst_2081 (
  .O(mux_o_2081),
  .I0(mux_o_1758),
  .I1(mux_o_1759),
  .S0(ad[5])
);
MUX2 mux_inst_2082 (
  .O(mux_o_2082),
  .I0(mux_o_1760),
  .I1(mux_o_1761),
  .S0(ad[5])
);
MUX2 mux_inst_2083 (
  .O(mux_o_2083),
  .I0(mux_o_1762),
  .I1(mux_o_1763),
  .S0(ad[5])
);
MUX2 mux_inst_2084 (
  .O(mux_o_2084),
  .I0(mux_o_1764),
  .I1(mux_o_1765),
  .S0(ad[5])
);
MUX2 mux_inst_2085 (
  .O(mux_o_2085),
  .I0(mux_o_1766),
  .I1(mux_o_1767),
  .S0(ad[5])
);
MUX2 mux_inst_2086 (
  .O(mux_o_2086),
  .I0(mux_o_1768),
  .I1(mux_o_1769),
  .S0(ad[5])
);
MUX2 mux_inst_2087 (
  .O(mux_o_2087),
  .I0(mux_o_1770),
  .I1(mux_o_1771),
  .S0(ad[5])
);
MUX2 mux_inst_2088 (
  .O(mux_o_2088),
  .I0(mux_o_1772),
  .I1(mux_o_1773),
  .S0(ad[5])
);
MUX2 mux_inst_2089 (
  .O(mux_o_2089),
  .I0(mux_o_1774),
  .I1(mux_o_1775),
  .S0(ad[5])
);
MUX2 mux_inst_2090 (
  .O(mux_o_2090),
  .I0(mux_o_1776),
  .I1(mux_o_1777),
  .S0(ad[5])
);
MUX2 mux_inst_2091 (
  .O(mux_o_2091),
  .I0(mux_o_1778),
  .I1(mux_o_1779),
  .S0(ad[5])
);
MUX2 mux_inst_2092 (
  .O(mux_o_2092),
  .I0(mux_o_1780),
  .I1(mux_o_1781),
  .S0(ad[5])
);
MUX2 mux_inst_2093 (
  .O(mux_o_2093),
  .I0(mux_o_1782),
  .I1(mux_o_1783),
  .S0(ad[5])
);
MUX2 mux_inst_2094 (
  .O(mux_o_2094),
  .I0(mux_o_1784),
  .I1(mux_o_1785),
  .S0(ad[5])
);
MUX2 mux_inst_2095 (
  .O(mux_o_2095),
  .I0(mux_o_1786),
  .I1(mux_o_1787),
  .S0(ad[5])
);
MUX2 mux_inst_2096 (
  .O(mux_o_2096),
  .I0(mux_o_1788),
  .I1(mux_o_1789),
  .S0(ad[5])
);
MUX2 mux_inst_2097 (
  .O(mux_o_2097),
  .I0(mux_o_1790),
  .I1(mux_o_1791),
  .S0(ad[5])
);
MUX2 mux_inst_2098 (
  .O(mux_o_2098),
  .I0(mux_o_1792),
  .I1(mux_o_1793),
  .S0(ad[5])
);
MUX2 mux_inst_2099 (
  .O(mux_o_2099),
  .I0(mux_o_1794),
  .I1(mux_o_1795),
  .S0(ad[5])
);
MUX2 mux_inst_2100 (
  .O(mux_o_2100),
  .I0(mux_o_1796),
  .I1(mux_o_1797),
  .S0(ad[5])
);
MUX2 mux_inst_2101 (
  .O(mux_o_2101),
  .I0(mux_o_1798),
  .I1(mux_o_1799),
  .S0(ad[5])
);
MUX2 mux_inst_2102 (
  .O(mux_o_2102),
  .I0(mux_o_1800),
  .I1(mux_o_1801),
  .S0(ad[5])
);
MUX2 mux_inst_2103 (
  .O(mux_o_2103),
  .I0(mux_o_1802),
  .I1(mux_o_1803),
  .S0(ad[5])
);
MUX2 mux_inst_2104 (
  .O(mux_o_2104),
  .I0(mux_o_1804),
  .I1(mux_o_1805),
  .S0(ad[5])
);
MUX2 mux_inst_2105 (
  .O(mux_o_2105),
  .I0(mux_o_1806),
  .I1(mux_o_1807),
  .S0(ad[5])
);
MUX2 mux_inst_2106 (
  .O(mux_o_2106),
  .I0(mux_o_1808),
  .I1(mux_o_1809),
  .S0(ad[5])
);
MUX2 mux_inst_2107 (
  .O(mux_o_2107),
  .I0(mux_o_1810),
  .I1(mux_o_1811),
  .S0(ad[5])
);
MUX2 mux_inst_2108 (
  .O(mux_o_2108),
  .I0(mux_o_1812),
  .I1(mux_o_1813),
  .S0(ad[5])
);
MUX2 mux_inst_2109 (
  .O(mux_o_2109),
  .I0(mux_o_1814),
  .I1(mux_o_1815),
  .S0(ad[5])
);
MUX2 mux_inst_2110 (
  .O(mux_o_2110),
  .I0(mux_o_1816),
  .I1(mux_o_1817),
  .S0(ad[5])
);
MUX2 mux_inst_2111 (
  .O(mux_o_2111),
  .I0(mux_o_1818),
  .I1(mux_o_1819),
  .S0(ad[5])
);
MUX2 mux_inst_2112 (
  .O(mux_o_2112),
  .I0(mux_o_1820),
  .I1(mux_o_1821),
  .S0(ad[5])
);
MUX2 mux_inst_2113 (
  .O(mux_o_2113),
  .I0(mux_o_1822),
  .I1(mux_o_1823),
  .S0(ad[5])
);
MUX2 mux_inst_2114 (
  .O(mux_o_2114),
  .I0(mux_o_1824),
  .I1(mux_o_1825),
  .S0(ad[5])
);
MUX2 mux_inst_2115 (
  .O(mux_o_2115),
  .I0(mux_o_1826),
  .I1(mux_o_1827),
  .S0(ad[5])
);
MUX2 mux_inst_2116 (
  .O(mux_o_2116),
  .I0(mux_o_1828),
  .I1(mux_o_1829),
  .S0(ad[5])
);
MUX2 mux_inst_2117 (
  .O(mux_o_2117),
  .I0(mux_o_1830),
  .I1(mux_o_1831),
  .S0(ad[5])
);
MUX2 mux_inst_2118 (
  .O(mux_o_2118),
  .I0(mux_o_1832),
  .I1(mux_o_1833),
  .S0(ad[5])
);
MUX2 mux_inst_2119 (
  .O(mux_o_2119),
  .I0(mux_o_1834),
  .I1(mux_o_1835),
  .S0(ad[5])
);
MUX2 mux_inst_2120 (
  .O(mux_o_2120),
  .I0(mux_o_1836),
  .I1(mux_o_1837),
  .S0(ad[5])
);
MUX2 mux_inst_2121 (
  .O(mux_o_2121),
  .I0(mux_o_1838),
  .I1(mux_o_1839),
  .S0(ad[5])
);
MUX2 mux_inst_2122 (
  .O(mux_o_2122),
  .I0(mux_o_1840),
  .I1(mux_o_1841),
  .S0(ad[5])
);
MUX2 mux_inst_2123 (
  .O(mux_o_2123),
  .I0(mux_o_1842),
  .I1(mux_o_1843),
  .S0(ad[5])
);
MUX2 mux_inst_2124 (
  .O(mux_o_2124),
  .I0(mux_o_1844),
  .I1(mux_o_1845),
  .S0(ad[5])
);
MUX2 mux_inst_2125 (
  .O(mux_o_2125),
  .I0(mux_o_1846),
  .I1(mux_o_1847),
  .S0(ad[5])
);
MUX2 mux_inst_2126 (
  .O(mux_o_2126),
  .I0(mux_o_1848),
  .I1(mux_o_1849),
  .S0(ad[5])
);
MUX2 mux_inst_2127 (
  .O(mux_o_2127),
  .I0(mux_o_1850),
  .I1(mux_o_1851),
  .S0(ad[5])
);
MUX2 mux_inst_2128 (
  .O(mux_o_2128),
  .I0(mux_o_1852),
  .I1(mux_o_1853),
  .S0(ad[5])
);
MUX2 mux_inst_2129 (
  .O(mux_o_2129),
  .I0(mux_o_1854),
  .I1(mux_o_1855),
  .S0(ad[5])
);
MUX2 mux_inst_2130 (
  .O(mux_o_2130),
  .I0(mux_o_1856),
  .I1(mux_o_1857),
  .S0(ad[5])
);
MUX2 mux_inst_2131 (
  .O(mux_o_2131),
  .I0(mux_o_1858),
  .I1(mux_o_1859),
  .S0(ad[5])
);
MUX2 mux_inst_2132 (
  .O(mux_o_2132),
  .I0(mux_o_1860),
  .I1(mux_o_1861),
  .S0(ad[5])
);
MUX2 mux_inst_2133 (
  .O(mux_o_2133),
  .I0(mux_o_1862),
  .I1(mux_o_1863),
  .S0(ad[5])
);
MUX2 mux_inst_2134 (
  .O(mux_o_2134),
  .I0(mux_o_1864),
  .I1(mux_o_1865),
  .S0(ad[5])
);
MUX2 mux_inst_2135 (
  .O(mux_o_2135),
  .I0(mux_o_1866),
  .I1(mux_o_1867),
  .S0(ad[5])
);
MUX2 mux_inst_2136 (
  .O(mux_o_2136),
  .I0(mux_o_1868),
  .I1(mux_o_1869),
  .S0(ad[5])
);
MUX2 mux_inst_2137 (
  .O(mux_o_2137),
  .I0(mux_o_1870),
  .I1(mux_o_1871),
  .S0(ad[5])
);
MUX2 mux_inst_2138 (
  .O(mux_o_2138),
  .I0(mux_o_1872),
  .I1(mux_o_1873),
  .S0(ad[5])
);
MUX2 mux_inst_2139 (
  .O(mux_o_2139),
  .I0(mux_o_1874),
  .I1(mux_o_1875),
  .S0(ad[5])
);
MUX2 mux_inst_2140 (
  .O(mux_o_2140),
  .I0(mux_o_1876),
  .I1(mux_o_1877),
  .S0(ad[5])
);
MUX2 mux_inst_2141 (
  .O(mux_o_2141),
  .I0(mux_o_1878),
  .I1(mux_o_1879),
  .S0(ad[5])
);
MUX2 mux_inst_2142 (
  .O(mux_o_2142),
  .I0(mux_o_1880),
  .I1(mux_o_1881),
  .S0(ad[5])
);
MUX2 mux_inst_2143 (
  .O(mux_o_2143),
  .I0(mux_o_1882),
  .I1(mux_o_1883),
  .S0(ad[5])
);
MUX2 mux_inst_2144 (
  .O(mux_o_2144),
  .I0(mux_o_1884),
  .I1(mux_o_1885),
  .S0(ad[5])
);
MUX2 mux_inst_2145 (
  .O(mux_o_2145),
  .I0(mux_o_1886),
  .I1(mux_o_1887),
  .S0(ad[5])
);
MUX2 mux_inst_2146 (
  .O(mux_o_2146),
  .I0(mux_o_1888),
  .I1(mux_o_1889),
  .S0(ad[5])
);
MUX2 mux_inst_2147 (
  .O(mux_o_2147),
  .I0(mux_o_1890),
  .I1(mux_o_1891),
  .S0(ad[5])
);
MUX2 mux_inst_2148 (
  .O(mux_o_2148),
  .I0(mux_o_1892),
  .I1(mux_o_1893),
  .S0(ad[5])
);
MUX2 mux_inst_2149 (
  .O(mux_o_2149),
  .I0(mux_o_1894),
  .I1(mux_o_1895),
  .S0(ad[5])
);
MUX2 mux_inst_2150 (
  .O(mux_o_2150),
  .I0(mux_o_1896),
  .I1(mux_o_1897),
  .S0(ad[5])
);
MUX2 mux_inst_2151 (
  .O(mux_o_2151),
  .I0(mux_o_1898),
  .I1(mux_o_1899),
  .S0(ad[5])
);
MUX2 mux_inst_2152 (
  .O(mux_o_2152),
  .I0(mux_o_1900),
  .I1(mux_o_1901),
  .S0(ad[5])
);
MUX2 mux_inst_2153 (
  .O(mux_o_2153),
  .I0(mux_o_1902),
  .I1(mux_o_1903),
  .S0(ad[5])
);
MUX2 mux_inst_2154 (
  .O(mux_o_2154),
  .I0(mux_o_1904),
  .I1(mux_o_1905),
  .S0(ad[5])
);
MUX2 mux_inst_2155 (
  .O(mux_o_2155),
  .I0(mux_o_1906),
  .I1(mux_o_1907),
  .S0(ad[5])
);
MUX2 mux_inst_2156 (
  .O(mux_o_2156),
  .I0(mux_o_1908),
  .I1(mux_o_1909),
  .S0(ad[5])
);
MUX2 mux_inst_2157 (
  .O(mux_o_2157),
  .I0(mux_o_1910),
  .I1(mux_o_1911),
  .S0(ad[5])
);
MUX2 mux_inst_2158 (
  .O(mux_o_2158),
  .I0(mux_o_1912),
  .I1(mux_o_1913),
  .S0(ad[5])
);
MUX2 mux_inst_2159 (
  .O(mux_o_2159),
  .I0(mux_o_1914),
  .I1(mux_o_1915),
  .S0(ad[5])
);
MUX2 mux_inst_2160 (
  .O(mux_o_2160),
  .I0(mux_o_1916),
  .I1(mux_o_1917),
  .S0(ad[5])
);
MUX2 mux_inst_2161 (
  .O(mux_o_2161),
  .I0(mux_o_1918),
  .I1(mux_o_1919),
  .S0(ad[5])
);
MUX2 mux_inst_2162 (
  .O(mux_o_2162),
  .I0(mux_o_1920),
  .I1(mux_o_1921),
  .S0(ad[5])
);
MUX2 mux_inst_2163 (
  .O(mux_o_2163),
  .I0(mux_o_1922),
  .I1(mux_o_1923),
  .S0(ad[5])
);
MUX2 mux_inst_2164 (
  .O(mux_o_2164),
  .I0(mux_o_1924),
  .I1(mux_o_1925),
  .S0(ad[5])
);
MUX2 mux_inst_2165 (
  .O(mux_o_2165),
  .I0(mux_o_1926),
  .I1(mux_o_1927),
  .S0(ad[5])
);
MUX2 mux_inst_2166 (
  .O(mux_o_2166),
  .I0(mux_o_1928),
  .I1(mux_o_1929),
  .S0(ad[5])
);
MUX2 mux_inst_2167 (
  .O(mux_o_2167),
  .I0(mux_o_1930),
  .I1(mux_o_1931),
  .S0(ad[5])
);
MUX2 mux_inst_2168 (
  .O(mux_o_2168),
  .I0(mux_o_1932),
  .I1(mux_o_1933),
  .S0(ad[5])
);
MUX2 mux_inst_2169 (
  .O(mux_o_2169),
  .I0(mux_o_1934),
  .I1(mux_o_1935),
  .S0(ad[5])
);
MUX2 mux_inst_2170 (
  .O(mux_o_2170),
  .I0(mux_o_1936),
  .I1(mux_o_1937),
  .S0(ad[5])
);
MUX2 mux_inst_2171 (
  .O(mux_o_2171),
  .I0(mux_o_1938),
  .I1(mux_o_1939),
  .S0(ad[5])
);
MUX2 mux_inst_2172 (
  .O(mux_o_2172),
  .I0(mux_o_1940),
  .I1(mux_o_1941),
  .S0(ad[5])
);
MUX2 mux_inst_2173 (
  .O(mux_o_2173),
  .I0(mux_o_1942),
  .I1(mux_o_1943),
  .S0(ad[5])
);
MUX2 mux_inst_2174 (
  .O(mux_o_2174),
  .I0(mux_o_1944),
  .I1(mux_o_1945),
  .S0(ad[5])
);
MUX2 mux_inst_2175 (
  .O(mux_o_2175),
  .I0(mux_o_1946),
  .I1(mux_o_1947),
  .S0(ad[5])
);
MUX2 mux_inst_2176 (
  .O(mux_o_2176),
  .I0(mux_o_1948),
  .I1(mux_o_1949),
  .S0(ad[5])
);
MUX2 mux_inst_2177 (
  .O(mux_o_2177),
  .I0(mux_o_1950),
  .I1(mux_o_1951),
  .S0(ad[5])
);
MUX2 mux_inst_2178 (
  .O(mux_o_2178),
  .I0(mux_o_1952),
  .I1(mux_o_1953),
  .S0(ad[5])
);
MUX2 mux_inst_2179 (
  .O(mux_o_2179),
  .I0(mux_o_1954),
  .I1(mux_o_1955),
  .S0(ad[5])
);
MUX2 mux_inst_2180 (
  .O(mux_o_2180),
  .I0(mux_o_1956),
  .I1(mux_o_1957),
  .S0(ad[5])
);
MUX2 mux_inst_2181 (
  .O(mux_o_2181),
  .I0(mux_o_1958),
  .I1(mux_o_1959),
  .S0(ad[5])
);
MUX2 mux_inst_2182 (
  .O(mux_o_2182),
  .I0(mux_o_1960),
  .I1(mux_o_1961),
  .S0(ad[5])
);
MUX2 mux_inst_2183 (
  .O(mux_o_2183),
  .I0(mux_o_1962),
  .I1(mux_o_1963),
  .S0(ad[5])
);
MUX2 mux_inst_2184 (
  .O(mux_o_2184),
  .I0(mux_o_1964),
  .I1(mux_o_1965),
  .S0(ad[5])
);
MUX2 mux_inst_2185 (
  .O(mux_o_2185),
  .I0(mux_o_1966),
  .I1(mux_o_1967),
  .S0(ad[5])
);
MUX2 mux_inst_2186 (
  .O(mux_o_2186),
  .I0(mux_o_1968),
  .I1(mux_o_1969),
  .S0(ad[5])
);
MUX2 mux_inst_2187 (
  .O(mux_o_2187),
  .I0(mux_o_1970),
  .I1(mux_o_1971),
  .S0(ad[5])
);
MUX2 mux_inst_2188 (
  .O(mux_o_2188),
  .I0(mux_o_1972),
  .I1(mux_o_1973),
  .S0(ad[5])
);
MUX2 mux_inst_2189 (
  .O(mux_o_2189),
  .I0(mux_o_1974),
  .I1(mux_o_1975),
  .S0(ad[5])
);
MUX2 mux_inst_2190 (
  .O(mux_o_2190),
  .I0(mux_o_1976),
  .I1(mux_o_1977),
  .S0(ad[5])
);
MUX2 mux_inst_2191 (
  .O(mux_o_2191),
  .I0(mux_o_1978),
  .I1(mux_o_1979),
  .S0(ad[5])
);
MUX2 mux_inst_2192 (
  .O(mux_o_2192),
  .I0(mux_o_1980),
  .I1(mux_o_1981),
  .S0(ad[5])
);
MUX2 mux_inst_2193 (
  .O(mux_o_2193),
  .I0(mux_o_1982),
  .I1(mux_o_1983),
  .S0(ad[5])
);
MUX2 mux_inst_2194 (
  .O(mux_o_2194),
  .I0(mux_o_1984),
  .I1(mux_o_1985),
  .S0(ad[5])
);
MUX2 mux_inst_2195 (
  .O(mux_o_2195),
  .I0(mux_o_1986),
  .I1(mux_o_1987),
  .S0(ad[5])
);
MUX2 mux_inst_2196 (
  .O(mux_o_2196),
  .I0(mux_o_1988),
  .I1(mux_o_1989),
  .S0(ad[5])
);
MUX2 mux_inst_2197 (
  .O(mux_o_2197),
  .I0(mux_o_1990),
  .I1(mux_o_1991),
  .S0(ad[5])
);
MUX2 mux_inst_2198 (
  .O(mux_o_2198),
  .I0(mux_o_1992),
  .I1(mux_o_1993),
  .S0(ad[5])
);
MUX2 mux_inst_2199 (
  .O(mux_o_2199),
  .I0(mux_o_1994),
  .I1(mux_o_1995),
  .S0(ad[5])
);
MUX2 mux_inst_2200 (
  .O(mux_o_2200),
  .I0(mux_o_1996),
  .I1(mux_o_1997),
  .S0(ad[5])
);
MUX2 mux_inst_2201 (
  .O(mux_o_2201),
  .I0(mux_o_1998),
  .I1(mux_o_1999),
  .S0(ad[5])
);
MUX2 mux_inst_2202 (
  .O(mux_o_2202),
  .I0(mux_o_2000),
  .I1(mux_o_2001),
  .S0(ad[5])
);
MUX2 mux_inst_2203 (
  .O(mux_o_2203),
  .I0(mux_o_2002),
  .I1(mux_o_2003),
  .S0(ad[5])
);
MUX2 mux_inst_2204 (
  .O(mux_o_2204),
  .I0(mux_o_2004),
  .I1(mux_o_2005),
  .S0(ad[6])
);
MUX2 mux_inst_2205 (
  .O(mux_o_2205),
  .I0(mux_o_2006),
  .I1(mux_o_2007),
  .S0(ad[6])
);
MUX2 mux_inst_2206 (
  .O(mux_o_2206),
  .I0(mux_o_2008),
  .I1(mux_o_2009),
  .S0(ad[6])
);
MUX2 mux_inst_2207 (
  .O(mux_o_2207),
  .I0(mux_o_2010),
  .I1(mux_o_2011),
  .S0(ad[6])
);
MUX2 mux_inst_2208 (
  .O(mux_o_2208),
  .I0(mux_o_2012),
  .I1(mux_o_2013),
  .S0(ad[6])
);
MUX2 mux_inst_2209 (
  .O(mux_o_2209),
  .I0(mux_o_2014),
  .I1(mux_o_2015),
  .S0(ad[6])
);
MUX2 mux_inst_2210 (
  .O(mux_o_2210),
  .I0(mux_o_2016),
  .I1(mux_o_2017),
  .S0(ad[6])
);
MUX2 mux_inst_2211 (
  .O(mux_o_2211),
  .I0(mux_o_2018),
  .I1(mux_o_2019),
  .S0(ad[6])
);
MUX2 mux_inst_2212 (
  .O(mux_o_2212),
  .I0(mux_o_2020),
  .I1(mux_o_2021),
  .S0(ad[6])
);
MUX2 mux_inst_2213 (
  .O(mux_o_2213),
  .I0(mux_o_2022),
  .I1(mux_o_2023),
  .S0(ad[6])
);
MUX2 mux_inst_2214 (
  .O(mux_o_2214),
  .I0(mux_o_2024),
  .I1(mux_o_2025),
  .S0(ad[6])
);
MUX2 mux_inst_2215 (
  .O(mux_o_2215),
  .I0(mux_o_2026),
  .I1(mux_o_2027),
  .S0(ad[6])
);
MUX2 mux_inst_2216 (
  .O(mux_o_2216),
  .I0(mux_o_2028),
  .I1(mux_o_2029),
  .S0(ad[6])
);
MUX2 mux_inst_2217 (
  .O(mux_o_2217),
  .I0(mux_o_2030),
  .I1(mux_o_2031),
  .S0(ad[6])
);
MUX2 mux_inst_2218 (
  .O(mux_o_2218),
  .I0(mux_o_2032),
  .I1(mux_o_2033),
  .S0(ad[6])
);
MUX2 mux_inst_2219 (
  .O(mux_o_2219),
  .I0(mux_o_2034),
  .I1(mux_o_2035),
  .S0(ad[6])
);
MUX2 mux_inst_2220 (
  .O(mux_o_2220),
  .I0(mux_o_2036),
  .I1(mux_o_2037),
  .S0(ad[6])
);
MUX2 mux_inst_2221 (
  .O(mux_o_2221),
  .I0(mux_o_2038),
  .I1(mux_o_2039),
  .S0(ad[6])
);
MUX2 mux_inst_2222 (
  .O(mux_o_2222),
  .I0(mux_o_2040),
  .I1(mux_o_2041),
  .S0(ad[6])
);
MUX2 mux_inst_2223 (
  .O(mux_o_2223),
  .I0(mux_o_2042),
  .I1(mux_o_2043),
  .S0(ad[6])
);
MUX2 mux_inst_2224 (
  .O(mux_o_2224),
  .I0(mux_o_2044),
  .I1(mux_o_2045),
  .S0(ad[6])
);
MUX2 mux_inst_2225 (
  .O(mux_o_2225),
  .I0(mux_o_2046),
  .I1(mux_o_2047),
  .S0(ad[6])
);
MUX2 mux_inst_2226 (
  .O(mux_o_2226),
  .I0(mux_o_2048),
  .I1(mux_o_2049),
  .S0(ad[6])
);
MUX2 mux_inst_2227 (
  .O(mux_o_2227),
  .I0(mux_o_2050),
  .I1(mux_o_2051),
  .S0(ad[6])
);
MUX2 mux_inst_2228 (
  .O(mux_o_2228),
  .I0(mux_o_2052),
  .I1(mux_o_2053),
  .S0(ad[6])
);
MUX2 mux_inst_2229 (
  .O(mux_o_2229),
  .I0(mux_o_2054),
  .I1(mux_o_2055),
  .S0(ad[6])
);
MUX2 mux_inst_2230 (
  .O(mux_o_2230),
  .I0(mux_o_2056),
  .I1(mux_o_2057),
  .S0(ad[6])
);
MUX2 mux_inst_2231 (
  .O(mux_o_2231),
  .I0(mux_o_2058),
  .I1(mux_o_2059),
  .S0(ad[6])
);
MUX2 mux_inst_2232 (
  .O(mux_o_2232),
  .I0(mux_o_2060),
  .I1(mux_o_2061),
  .S0(ad[6])
);
MUX2 mux_inst_2233 (
  .O(mux_o_2233),
  .I0(mux_o_2062),
  .I1(mux_o_2063),
  .S0(ad[6])
);
MUX2 mux_inst_2234 (
  .O(mux_o_2234),
  .I0(mux_o_2064),
  .I1(mux_o_2065),
  .S0(ad[6])
);
MUX2 mux_inst_2235 (
  .O(mux_o_2235),
  .I0(mux_o_2066),
  .I1(mux_o_2067),
  .S0(ad[6])
);
MUX2 mux_inst_2236 (
  .O(mux_o_2236),
  .I0(mux_o_2068),
  .I1(mux_o_2069),
  .S0(ad[6])
);
MUX2 mux_inst_2237 (
  .O(mux_o_2237),
  .I0(mux_o_2070),
  .I1(mux_o_2071),
  .S0(ad[6])
);
MUX2 mux_inst_2238 (
  .O(mux_o_2238),
  .I0(mux_o_2072),
  .I1(mux_o_2073),
  .S0(ad[6])
);
MUX2 mux_inst_2239 (
  .O(mux_o_2239),
  .I0(mux_o_2074),
  .I1(mux_o_2075),
  .S0(ad[6])
);
MUX2 mux_inst_2240 (
  .O(mux_o_2240),
  .I0(mux_o_2076),
  .I1(mux_o_2077),
  .S0(ad[6])
);
MUX2 mux_inst_2241 (
  .O(mux_o_2241),
  .I0(mux_o_2078),
  .I1(mux_o_2079),
  .S0(ad[6])
);
MUX2 mux_inst_2242 (
  .O(mux_o_2242),
  .I0(mux_o_2080),
  .I1(mux_o_2081),
  .S0(ad[6])
);
MUX2 mux_inst_2243 (
  .O(mux_o_2243),
  .I0(mux_o_2082),
  .I1(mux_o_2083),
  .S0(ad[6])
);
MUX2 mux_inst_2244 (
  .O(mux_o_2244),
  .I0(mux_o_2084),
  .I1(mux_o_2085),
  .S0(ad[6])
);
MUX2 mux_inst_2245 (
  .O(mux_o_2245),
  .I0(mux_o_2086),
  .I1(mux_o_2087),
  .S0(ad[6])
);
MUX2 mux_inst_2246 (
  .O(mux_o_2246),
  .I0(mux_o_2088),
  .I1(mux_o_2089),
  .S0(ad[6])
);
MUX2 mux_inst_2247 (
  .O(mux_o_2247),
  .I0(mux_o_2090),
  .I1(mux_o_2091),
  .S0(ad[6])
);
MUX2 mux_inst_2248 (
  .O(mux_o_2248),
  .I0(mux_o_2092),
  .I1(mux_o_2093),
  .S0(ad[6])
);
MUX2 mux_inst_2249 (
  .O(mux_o_2249),
  .I0(mux_o_2094),
  .I1(mux_o_2095),
  .S0(ad[6])
);
MUX2 mux_inst_2250 (
  .O(mux_o_2250),
  .I0(mux_o_2096),
  .I1(mux_o_2097),
  .S0(ad[6])
);
MUX2 mux_inst_2251 (
  .O(mux_o_2251),
  .I0(mux_o_2098),
  .I1(mux_o_2099),
  .S0(ad[6])
);
MUX2 mux_inst_2252 (
  .O(mux_o_2252),
  .I0(mux_o_2100),
  .I1(mux_o_2101),
  .S0(ad[6])
);
MUX2 mux_inst_2253 (
  .O(mux_o_2253),
  .I0(mux_o_2102),
  .I1(mux_o_2103),
  .S0(ad[6])
);
MUX2 mux_inst_2254 (
  .O(mux_o_2254),
  .I0(mux_o_2104),
  .I1(mux_o_2105),
  .S0(ad[6])
);
MUX2 mux_inst_2255 (
  .O(mux_o_2255),
  .I0(mux_o_2106),
  .I1(mux_o_2107),
  .S0(ad[6])
);
MUX2 mux_inst_2256 (
  .O(mux_o_2256),
  .I0(mux_o_2108),
  .I1(mux_o_2109),
  .S0(ad[6])
);
MUX2 mux_inst_2257 (
  .O(mux_o_2257),
  .I0(mux_o_2110),
  .I1(mux_o_2111),
  .S0(ad[6])
);
MUX2 mux_inst_2258 (
  .O(mux_o_2258),
  .I0(mux_o_2112),
  .I1(mux_o_2113),
  .S0(ad[6])
);
MUX2 mux_inst_2259 (
  .O(mux_o_2259),
  .I0(mux_o_2114),
  .I1(mux_o_2115),
  .S0(ad[6])
);
MUX2 mux_inst_2260 (
  .O(mux_o_2260),
  .I0(mux_o_2116),
  .I1(mux_o_2117),
  .S0(ad[6])
);
MUX2 mux_inst_2261 (
  .O(mux_o_2261),
  .I0(mux_o_2118),
  .I1(mux_o_2119),
  .S0(ad[6])
);
MUX2 mux_inst_2262 (
  .O(mux_o_2262),
  .I0(mux_o_2120),
  .I1(mux_o_2121),
  .S0(ad[6])
);
MUX2 mux_inst_2263 (
  .O(mux_o_2263),
  .I0(mux_o_2122),
  .I1(mux_o_2123),
  .S0(ad[6])
);
MUX2 mux_inst_2264 (
  .O(mux_o_2264),
  .I0(mux_o_2124),
  .I1(mux_o_2125),
  .S0(ad[6])
);
MUX2 mux_inst_2265 (
  .O(mux_o_2265),
  .I0(mux_o_2126),
  .I1(mux_o_2127),
  .S0(ad[6])
);
MUX2 mux_inst_2266 (
  .O(mux_o_2266),
  .I0(mux_o_2128),
  .I1(mux_o_2129),
  .S0(ad[6])
);
MUX2 mux_inst_2267 (
  .O(mux_o_2267),
  .I0(mux_o_2130),
  .I1(mux_o_2131),
  .S0(ad[6])
);
MUX2 mux_inst_2268 (
  .O(mux_o_2268),
  .I0(mux_o_2132),
  .I1(mux_o_2133),
  .S0(ad[6])
);
MUX2 mux_inst_2269 (
  .O(mux_o_2269),
  .I0(mux_o_2134),
  .I1(mux_o_2135),
  .S0(ad[6])
);
MUX2 mux_inst_2270 (
  .O(mux_o_2270),
  .I0(mux_o_2136),
  .I1(mux_o_2137),
  .S0(ad[6])
);
MUX2 mux_inst_2271 (
  .O(mux_o_2271),
  .I0(mux_o_2138),
  .I1(mux_o_2139),
  .S0(ad[6])
);
MUX2 mux_inst_2272 (
  .O(mux_o_2272),
  .I0(mux_o_2140),
  .I1(mux_o_2141),
  .S0(ad[6])
);
MUX2 mux_inst_2273 (
  .O(mux_o_2273),
  .I0(mux_o_2142),
  .I1(mux_o_2143),
  .S0(ad[6])
);
MUX2 mux_inst_2274 (
  .O(mux_o_2274),
  .I0(mux_o_2144),
  .I1(mux_o_2145),
  .S0(ad[6])
);
MUX2 mux_inst_2275 (
  .O(mux_o_2275),
  .I0(mux_o_2146),
  .I1(mux_o_2147),
  .S0(ad[6])
);
MUX2 mux_inst_2276 (
  .O(mux_o_2276),
  .I0(mux_o_2148),
  .I1(mux_o_2149),
  .S0(ad[6])
);
MUX2 mux_inst_2277 (
  .O(mux_o_2277),
  .I0(mux_o_2150),
  .I1(mux_o_2151),
  .S0(ad[6])
);
MUX2 mux_inst_2278 (
  .O(mux_o_2278),
  .I0(mux_o_2152),
  .I1(mux_o_2153),
  .S0(ad[6])
);
MUX2 mux_inst_2279 (
  .O(mux_o_2279),
  .I0(mux_o_2154),
  .I1(mux_o_2155),
  .S0(ad[6])
);
MUX2 mux_inst_2280 (
  .O(mux_o_2280),
  .I0(mux_o_2156),
  .I1(mux_o_2157),
  .S0(ad[6])
);
MUX2 mux_inst_2281 (
  .O(mux_o_2281),
  .I0(mux_o_2158),
  .I1(mux_o_2159),
  .S0(ad[6])
);
MUX2 mux_inst_2282 (
  .O(mux_o_2282),
  .I0(mux_o_2160),
  .I1(mux_o_2161),
  .S0(ad[6])
);
MUX2 mux_inst_2283 (
  .O(mux_o_2283),
  .I0(mux_o_2162),
  .I1(mux_o_2163),
  .S0(ad[6])
);
MUX2 mux_inst_2284 (
  .O(mux_o_2284),
  .I0(mux_o_2164),
  .I1(mux_o_2165),
  .S0(ad[6])
);
MUX2 mux_inst_2285 (
  .O(mux_o_2285),
  .I0(mux_o_2166),
  .I1(mux_o_2167),
  .S0(ad[6])
);
MUX2 mux_inst_2286 (
  .O(mux_o_2286),
  .I0(mux_o_2168),
  .I1(mux_o_2169),
  .S0(ad[6])
);
MUX2 mux_inst_2287 (
  .O(mux_o_2287),
  .I0(mux_o_2170),
  .I1(mux_o_2171),
  .S0(ad[6])
);
MUX2 mux_inst_2288 (
  .O(mux_o_2288),
  .I0(mux_o_2172),
  .I1(mux_o_2173),
  .S0(ad[6])
);
MUX2 mux_inst_2289 (
  .O(mux_o_2289),
  .I0(mux_o_2174),
  .I1(mux_o_2175),
  .S0(ad[6])
);
MUX2 mux_inst_2290 (
  .O(mux_o_2290),
  .I0(mux_o_2176),
  .I1(mux_o_2177),
  .S0(ad[6])
);
MUX2 mux_inst_2291 (
  .O(mux_o_2291),
  .I0(mux_o_2178),
  .I1(mux_o_2179),
  .S0(ad[6])
);
MUX2 mux_inst_2292 (
  .O(mux_o_2292),
  .I0(mux_o_2180),
  .I1(mux_o_2181),
  .S0(ad[6])
);
MUX2 mux_inst_2293 (
  .O(mux_o_2293),
  .I0(mux_o_2182),
  .I1(mux_o_2183),
  .S0(ad[6])
);
MUX2 mux_inst_2294 (
  .O(mux_o_2294),
  .I0(mux_o_2184),
  .I1(mux_o_2185),
  .S0(ad[6])
);
MUX2 mux_inst_2295 (
  .O(mux_o_2295),
  .I0(mux_o_2186),
  .I1(mux_o_2187),
  .S0(ad[6])
);
MUX2 mux_inst_2296 (
  .O(mux_o_2296),
  .I0(mux_o_2188),
  .I1(mux_o_2189),
  .S0(ad[6])
);
MUX2 mux_inst_2297 (
  .O(mux_o_2297),
  .I0(mux_o_2190),
  .I1(mux_o_2191),
  .S0(ad[6])
);
MUX2 mux_inst_2298 (
  .O(mux_o_2298),
  .I0(mux_o_2192),
  .I1(mux_o_2193),
  .S0(ad[6])
);
MUX2 mux_inst_2299 (
  .O(mux_o_2299),
  .I0(mux_o_2194),
  .I1(mux_o_2195),
  .S0(ad[6])
);
MUX2 mux_inst_2300 (
  .O(mux_o_2300),
  .I0(mux_o_2196),
  .I1(mux_o_2197),
  .S0(ad[6])
);
MUX2 mux_inst_2301 (
  .O(mux_o_2301),
  .I0(mux_o_2198),
  .I1(mux_o_2199),
  .S0(ad[6])
);
MUX2 mux_inst_2302 (
  .O(mux_o_2302),
  .I0(mux_o_2200),
  .I1(mux_o_2201),
  .S0(ad[6])
);
MUX2 mux_inst_2303 (
  .O(mux_o_2303),
  .I0(mux_o_2202),
  .I1(mux_o_2203),
  .S0(ad[6])
);
MUX2 mux_inst_2304 (
  .O(mux_o_2304),
  .I0(mux_o_2204),
  .I1(mux_o_2205),
  .S0(ad[7])
);
MUX2 mux_inst_2305 (
  .O(mux_o_2305),
  .I0(mux_o_2206),
  .I1(mux_o_2207),
  .S0(ad[7])
);
MUX2 mux_inst_2306 (
  .O(mux_o_2306),
  .I0(mux_o_2208),
  .I1(mux_o_2209),
  .S0(ad[7])
);
MUX2 mux_inst_2307 (
  .O(mux_o_2307),
  .I0(mux_o_2210),
  .I1(mux_o_2211),
  .S0(ad[7])
);
MUX2 mux_inst_2308 (
  .O(mux_o_2308),
  .I0(mux_o_2212),
  .I1(mux_o_2213),
  .S0(ad[7])
);
MUX2 mux_inst_2309 (
  .O(mux_o_2309),
  .I0(mux_o_2214),
  .I1(mux_o_2215),
  .S0(ad[7])
);
MUX2 mux_inst_2310 (
  .O(mux_o_2310),
  .I0(mux_o_2216),
  .I1(mux_o_2217),
  .S0(ad[7])
);
MUX2 mux_inst_2311 (
  .O(mux_o_2311),
  .I0(mux_o_2218),
  .I1(mux_o_2219),
  .S0(ad[7])
);
MUX2 mux_inst_2312 (
  .O(mux_o_2312),
  .I0(mux_o_2220),
  .I1(mux_o_2221),
  .S0(ad[7])
);
MUX2 mux_inst_2313 (
  .O(mux_o_2313),
  .I0(mux_o_2222),
  .I1(mux_o_2223),
  .S0(ad[7])
);
MUX2 mux_inst_2314 (
  .O(mux_o_2314),
  .I0(mux_o_2224),
  .I1(mux_o_2225),
  .S0(ad[7])
);
MUX2 mux_inst_2315 (
  .O(mux_o_2315),
  .I0(mux_o_2226),
  .I1(mux_o_2227),
  .S0(ad[7])
);
MUX2 mux_inst_2316 (
  .O(mux_o_2316),
  .I0(mux_o_2228),
  .I1(mux_o_2229),
  .S0(ad[7])
);
MUX2 mux_inst_2317 (
  .O(mux_o_2317),
  .I0(mux_o_2230),
  .I1(mux_o_2231),
  .S0(ad[7])
);
MUX2 mux_inst_2318 (
  .O(mux_o_2318),
  .I0(mux_o_2232),
  .I1(mux_o_2233),
  .S0(ad[7])
);
MUX2 mux_inst_2319 (
  .O(mux_o_2319),
  .I0(mux_o_2234),
  .I1(mux_o_2235),
  .S0(ad[7])
);
MUX2 mux_inst_2320 (
  .O(mux_o_2320),
  .I0(mux_o_2236),
  .I1(mux_o_2237),
  .S0(ad[7])
);
MUX2 mux_inst_2321 (
  .O(mux_o_2321),
  .I0(mux_o_2238),
  .I1(mux_o_2239),
  .S0(ad[7])
);
MUX2 mux_inst_2322 (
  .O(mux_o_2322),
  .I0(mux_o_2240),
  .I1(mux_o_2241),
  .S0(ad[7])
);
MUX2 mux_inst_2323 (
  .O(mux_o_2323),
  .I0(mux_o_2242),
  .I1(mux_o_2243),
  .S0(ad[7])
);
MUX2 mux_inst_2324 (
  .O(mux_o_2324),
  .I0(mux_o_2244),
  .I1(mux_o_2245),
  .S0(ad[7])
);
MUX2 mux_inst_2325 (
  .O(mux_o_2325),
  .I0(mux_o_2246),
  .I1(mux_o_2247),
  .S0(ad[7])
);
MUX2 mux_inst_2326 (
  .O(mux_o_2326),
  .I0(mux_o_2248),
  .I1(mux_o_2249),
  .S0(ad[7])
);
MUX2 mux_inst_2327 (
  .O(mux_o_2327),
  .I0(mux_o_2250),
  .I1(mux_o_2251),
  .S0(ad[7])
);
MUX2 mux_inst_2328 (
  .O(mux_o_2328),
  .I0(mux_o_2252),
  .I1(mux_o_2253),
  .S0(ad[7])
);
MUX2 mux_inst_2329 (
  .O(mux_o_2329),
  .I0(mux_o_2254),
  .I1(mux_o_2255),
  .S0(ad[7])
);
MUX2 mux_inst_2330 (
  .O(mux_o_2330),
  .I0(mux_o_2256),
  .I1(mux_o_2257),
  .S0(ad[7])
);
MUX2 mux_inst_2331 (
  .O(mux_o_2331),
  .I0(mux_o_2258),
  .I1(mux_o_2259),
  .S0(ad[7])
);
MUX2 mux_inst_2332 (
  .O(mux_o_2332),
  .I0(mux_o_2260),
  .I1(mux_o_2261),
  .S0(ad[7])
);
MUX2 mux_inst_2333 (
  .O(mux_o_2333),
  .I0(mux_o_2262),
  .I1(mux_o_2263),
  .S0(ad[7])
);
MUX2 mux_inst_2334 (
  .O(mux_o_2334),
  .I0(mux_o_2264),
  .I1(mux_o_2265),
  .S0(ad[7])
);
MUX2 mux_inst_2335 (
  .O(mux_o_2335),
  .I0(mux_o_2266),
  .I1(mux_o_2267),
  .S0(ad[7])
);
MUX2 mux_inst_2336 (
  .O(mux_o_2336),
  .I0(mux_o_2268),
  .I1(mux_o_2269),
  .S0(ad[7])
);
MUX2 mux_inst_2337 (
  .O(mux_o_2337),
  .I0(mux_o_2270),
  .I1(mux_o_2271),
  .S0(ad[7])
);
MUX2 mux_inst_2338 (
  .O(mux_o_2338),
  .I0(mux_o_2272),
  .I1(mux_o_2273),
  .S0(ad[7])
);
MUX2 mux_inst_2339 (
  .O(mux_o_2339),
  .I0(mux_o_2274),
  .I1(mux_o_2275),
  .S0(ad[7])
);
MUX2 mux_inst_2340 (
  .O(mux_o_2340),
  .I0(mux_o_2276),
  .I1(mux_o_2277),
  .S0(ad[7])
);
MUX2 mux_inst_2341 (
  .O(mux_o_2341),
  .I0(mux_o_2278),
  .I1(mux_o_2279),
  .S0(ad[7])
);
MUX2 mux_inst_2342 (
  .O(mux_o_2342),
  .I0(mux_o_2280),
  .I1(mux_o_2281),
  .S0(ad[7])
);
MUX2 mux_inst_2343 (
  .O(mux_o_2343),
  .I0(mux_o_2282),
  .I1(mux_o_2283),
  .S0(ad[7])
);
MUX2 mux_inst_2344 (
  .O(mux_o_2344),
  .I0(mux_o_2284),
  .I1(mux_o_2285),
  .S0(ad[7])
);
MUX2 mux_inst_2345 (
  .O(mux_o_2345),
  .I0(mux_o_2286),
  .I1(mux_o_2287),
  .S0(ad[7])
);
MUX2 mux_inst_2346 (
  .O(mux_o_2346),
  .I0(mux_o_2288),
  .I1(mux_o_2289),
  .S0(ad[7])
);
MUX2 mux_inst_2347 (
  .O(mux_o_2347),
  .I0(mux_o_2290),
  .I1(mux_o_2291),
  .S0(ad[7])
);
MUX2 mux_inst_2348 (
  .O(mux_o_2348),
  .I0(mux_o_2292),
  .I1(mux_o_2293),
  .S0(ad[7])
);
MUX2 mux_inst_2349 (
  .O(mux_o_2349),
  .I0(mux_o_2294),
  .I1(mux_o_2295),
  .S0(ad[7])
);
MUX2 mux_inst_2350 (
  .O(mux_o_2350),
  .I0(mux_o_2296),
  .I1(mux_o_2297),
  .S0(ad[7])
);
MUX2 mux_inst_2351 (
  .O(mux_o_2351),
  .I0(mux_o_2298),
  .I1(mux_o_2299),
  .S0(ad[7])
);
MUX2 mux_inst_2352 (
  .O(mux_o_2352),
  .I0(mux_o_2300),
  .I1(mux_o_2301),
  .S0(ad[7])
);
MUX2 mux_inst_2353 (
  .O(mux_o_2353),
  .I0(mux_o_2302),
  .I1(mux_o_2303),
  .S0(ad[7])
);
MUX2 mux_inst_2354 (
  .O(mux_o_2354),
  .I0(mux_o_2304),
  .I1(mux_o_2305),
  .S0(ad[8])
);
MUX2 mux_inst_2355 (
  .O(mux_o_2355),
  .I0(mux_o_2306),
  .I1(mux_o_2307),
  .S0(ad[8])
);
MUX2 mux_inst_2356 (
  .O(mux_o_2356),
  .I0(mux_o_2308),
  .I1(mux_o_2309),
  .S0(ad[8])
);
MUX2 mux_inst_2357 (
  .O(mux_o_2357),
  .I0(mux_o_2310),
  .I1(mux_o_2311),
  .S0(ad[8])
);
MUX2 mux_inst_2358 (
  .O(mux_o_2358),
  .I0(mux_o_2312),
  .I1(mux_o_2313),
  .S0(ad[8])
);
MUX2 mux_inst_2359 (
  .O(mux_o_2359),
  .I0(mux_o_2314),
  .I1(mux_o_2315),
  .S0(ad[8])
);
MUX2 mux_inst_2360 (
  .O(mux_o_2360),
  .I0(mux_o_2316),
  .I1(mux_o_2317),
  .S0(ad[8])
);
MUX2 mux_inst_2361 (
  .O(mux_o_2361),
  .I0(mux_o_2318),
  .I1(mux_o_2319),
  .S0(ad[8])
);
MUX2 mux_inst_2362 (
  .O(mux_o_2362),
  .I0(mux_o_2320),
  .I1(mux_o_2321),
  .S0(ad[8])
);
MUX2 mux_inst_2363 (
  .O(mux_o_2363),
  .I0(mux_o_2322),
  .I1(mux_o_2323),
  .S0(ad[8])
);
MUX2 mux_inst_2364 (
  .O(mux_o_2364),
  .I0(mux_o_2324),
  .I1(mux_o_2325),
  .S0(ad[8])
);
MUX2 mux_inst_2365 (
  .O(mux_o_2365),
  .I0(mux_o_2326),
  .I1(mux_o_2327),
  .S0(ad[8])
);
MUX2 mux_inst_2366 (
  .O(mux_o_2366),
  .I0(mux_o_2328),
  .I1(mux_o_2329),
  .S0(ad[8])
);
MUX2 mux_inst_2367 (
  .O(mux_o_2367),
  .I0(mux_o_2330),
  .I1(mux_o_2331),
  .S0(ad[8])
);
MUX2 mux_inst_2368 (
  .O(mux_o_2368),
  .I0(mux_o_2332),
  .I1(mux_o_2333),
  .S0(ad[8])
);
MUX2 mux_inst_2369 (
  .O(mux_o_2369),
  .I0(mux_o_2334),
  .I1(mux_o_2335),
  .S0(ad[8])
);
MUX2 mux_inst_2370 (
  .O(mux_o_2370),
  .I0(mux_o_2336),
  .I1(mux_o_2337),
  .S0(ad[8])
);
MUX2 mux_inst_2371 (
  .O(mux_o_2371),
  .I0(mux_o_2338),
  .I1(mux_o_2339),
  .S0(ad[8])
);
MUX2 mux_inst_2372 (
  .O(mux_o_2372),
  .I0(mux_o_2340),
  .I1(mux_o_2341),
  .S0(ad[8])
);
MUX2 mux_inst_2373 (
  .O(mux_o_2373),
  .I0(mux_o_2342),
  .I1(mux_o_2343),
  .S0(ad[8])
);
MUX2 mux_inst_2374 (
  .O(mux_o_2374),
  .I0(mux_o_2344),
  .I1(mux_o_2345),
  .S0(ad[8])
);
MUX2 mux_inst_2375 (
  .O(mux_o_2375),
  .I0(mux_o_2346),
  .I1(mux_o_2347),
  .S0(ad[8])
);
MUX2 mux_inst_2376 (
  .O(mux_o_2376),
  .I0(mux_o_2348),
  .I1(mux_o_2349),
  .S0(ad[8])
);
MUX2 mux_inst_2377 (
  .O(mux_o_2377),
  .I0(mux_o_2350),
  .I1(mux_o_2351),
  .S0(ad[8])
);
MUX2 mux_inst_2378 (
  .O(mux_o_2378),
  .I0(mux_o_2352),
  .I1(mux_o_2353),
  .S0(ad[8])
);
MUX2 mux_inst_2379 (
  .O(mux_o_2379),
  .I0(mux_o_2354),
  .I1(mux_o_2355),
  .S0(ad[9])
);
MUX2 mux_inst_2380 (
  .O(mux_o_2380),
  .I0(mux_o_2356),
  .I1(mux_o_2357),
  .S0(ad[9])
);
MUX2 mux_inst_2381 (
  .O(mux_o_2381),
  .I0(mux_o_2358),
  .I1(mux_o_2359),
  .S0(ad[9])
);
MUX2 mux_inst_2382 (
  .O(mux_o_2382),
  .I0(mux_o_2360),
  .I1(mux_o_2361),
  .S0(ad[9])
);
MUX2 mux_inst_2383 (
  .O(mux_o_2383),
  .I0(mux_o_2362),
  .I1(mux_o_2363),
  .S0(ad[9])
);
MUX2 mux_inst_2384 (
  .O(mux_o_2384),
  .I0(mux_o_2364),
  .I1(mux_o_2365),
  .S0(ad[9])
);
MUX2 mux_inst_2385 (
  .O(mux_o_2385),
  .I0(mux_o_2366),
  .I1(mux_o_2367),
  .S0(ad[9])
);
MUX2 mux_inst_2386 (
  .O(mux_o_2386),
  .I0(mux_o_2368),
  .I1(mux_o_2369),
  .S0(ad[9])
);
MUX2 mux_inst_2387 (
  .O(mux_o_2387),
  .I0(mux_o_2370),
  .I1(mux_o_2371),
  .S0(ad[9])
);
MUX2 mux_inst_2388 (
  .O(mux_o_2388),
  .I0(mux_o_2372),
  .I1(mux_o_2373),
  .S0(ad[9])
);
MUX2 mux_inst_2389 (
  .O(mux_o_2389),
  .I0(mux_o_2374),
  .I1(mux_o_2375),
  .S0(ad[9])
);
MUX2 mux_inst_2390 (
  .O(mux_o_2390),
  .I0(mux_o_2376),
  .I1(mux_o_2377),
  .S0(ad[9])
);
MUX2 mux_inst_2392 (
  .O(mux_o_2392),
  .I0(mux_o_2379),
  .I1(mux_o_2380),
  .S0(ad[10])
);
MUX2 mux_inst_2393 (
  .O(mux_o_2393),
  .I0(mux_o_2381),
  .I1(mux_o_2382),
  .S0(ad[10])
);
MUX2 mux_inst_2394 (
  .O(mux_o_2394),
  .I0(mux_o_2383),
  .I1(mux_o_2384),
  .S0(ad[10])
);
MUX2 mux_inst_2395 (
  .O(mux_o_2395),
  .I0(mux_o_2385),
  .I1(mux_o_2386),
  .S0(ad[10])
);
MUX2 mux_inst_2396 (
  .O(mux_o_2396),
  .I0(mux_o_2387),
  .I1(mux_o_2388),
  .S0(ad[10])
);
MUX2 mux_inst_2397 (
  .O(mux_o_2397),
  .I0(mux_o_2389),
  .I1(mux_o_2390),
  .S0(ad[10])
);
MUX2 mux_inst_2399 (
  .O(mux_o_2399),
  .I0(mux_o_2392),
  .I1(mux_o_2393),
  .S0(ad[11])
);
MUX2 mux_inst_2400 (
  .O(mux_o_2400),
  .I0(mux_o_2394),
  .I1(mux_o_2395),
  .S0(ad[11])
);
MUX2 mux_inst_2401 (
  .O(mux_o_2401),
  .I0(mux_o_2396),
  .I1(mux_o_2397),
  .S0(ad[11])
);
MUX2 mux_inst_2403 (
  .O(mux_o_2403),
  .I0(mux_o_2399),
  .I1(mux_o_2400),
  .S0(ad[12])
);
MUX2 mux_inst_2404 (
  .O(mux_o_2404),
  .I0(mux_o_2401),
  .I1(mux_o_2378),
  .S0(ad[12])
);
MUX2 mux_inst_2405 (
  .O(dout[2]),
  .I0(mux_o_2403),
  .I1(mux_o_2404),
  .S0(ad[13])
);
endmodule //Gowin_RAM16S
